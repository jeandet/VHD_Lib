-- FillFifo.vhd
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FillFifo is
generic(
    Data_sz  : integer range 1 to 32 := 16;
    Fifo_cnt : integer range 1 to 8 := 5
    );
port(
    clk         : in std_logic;
    raz        : in std_logic;
    write : out std_logic_vector(Fifo_cnt-1 downto 0);
    reuse : out std_logic_vector(Fifo_cnt-1 downto 0);
    data : out std_logic_vector(Fifo_cnt*Data_sz-1 downto 0)
);
end entity;


architecture ar_FillFifo of FillFifo is

signal i : integer := 0;

type etat is (eX,e0,e00);
signal ect : etat;

type Tbl is array(natural range <>) of std_logic_vector(Data_sz-1 downto 0);

--constant TblA : Tbl (0 to 255) := (X"FFFF",X"0142",X"0282",X"03C2",X"04FF",X"0638",X"076E",X"08A0",X"09CC",X"0AF2",X"0C11",X"0D29",X"0E39",X"0F40",X"103E",X"1131",X"121A",X"12F8",X"13CA",X"1490",X"1549",X"15F5",X"1694",X"1724",X"17A7",X"181B",X"187F",X"18D5",X"191C",X"1953",X"197A",X"1992",X"199A",X"1992",X"197A",X"1953",X"191C",X"18D5",X"187F",X"181B",X"17A7",X"1724",X"1694",X"15F5",X"1549",X"1490",X"13CA",X"12F8",X"121A",X"1131",X"103E",X"0F40",X"0E39",X"0D29",X"0C11",X"0AF2",X"09CC",X"08A0",X"076E",X"0638",X"04FF",X"03C2",X"0282",X"0142",X"0000",X"FEBE",X"FD7E",X"FC3E",X"FB01",X"F9C8",X"F892",X"F760",X"F634",X"F50E",X"F3EF",X"F2D7",X"F1C7",X"F0C0",X"EFC2",X"EECF",X"EDE6",X"ED08",X"EC36",X"EB70",X"EAB7",X"EA0B",X"E96C",X"E8DC",X"E859",X"E7E5",X"E781",X"E72B",X"E6E4",X"E6AD",X"E686",X"E66E",X"E666",X"E66E",X"E686",X"E6AD",X"E6E4",X"E72B",X"E781",X"E7E5",X"E859",X"E8DC",X"E96C",X"EA0B",X"EAB7",X"EB70",X"EC36",X"ED08",X"EDE6",X"EECF",X"EFC2",X"F0C0",X"F1C7",X"F2D7",X"F3EF",X"F50E",X"F634",X"F760",X"F892",X"F9C8",X"FB01",X"FC3E",X"FD7E",X"FEBE",X"0000",X"0142",X"0282",X"03C2",X"04FF",X"0638",X"076E",X"08A0",X"09CC",X"0AF2",X"0C11",X"0D29",X"0E39",X"0F40",X"103E",X"1131",X"121A",X"12F8",X"13CA",X"1490",X"1549",X"15F5",X"1694",X"1724",X"17A7",X"181B",X"187F",X"18D5",X"191C",X"1953",X"197A",X"1992",X"199A",X"1992",X"197A",X"1953",X"191C",X"18D5",X"187F",X"181B",X"17A7",X"1724",X"1694",X"15F5",X"1549",X"1490",X"13CA",X"12F8",X"121A",X"1131",X"103E",X"0F40",X"0E39",X"0D29",X"0C11",X"0AF2",X"09CC",X"08A0",X"076E",X"0638",X"04FF",X"03C2",X"0282",X"0142",X"0000",X"FEBE",X"FD7E",X"FC3E",X"FB01",X"F9C8",X"F892",X"F760",X"F634",X"F50E",X"F3EF",X"F2D7",X"F1C7",X"F0C0",X"EFC2",X"EECF",X"EDE6",X"ED08",X"EC36",X"EB70",X"EAB7",X"EA0B",X"E96C",X"E8DC",X"E859",X"E7E5",X"E781",X"E72B", 
--X"E6E4",X"E6AD",X"E686",X"E66E",X"E666",X"E66E",X"E686",X"E6AD",X"E6E4",X"E72B",X"E781",X"E7E5",X"E859",X"E8DC",X"E96C",X"EA0B",X"EAB7",X"EB70",X"EC36",X"ED08",X"EDE6",X"EECF",X"EFC2",X"F0C0",X"F1C7",X"F2D7",X"F3EF",X"F50E",X"F634",X"F760",X"F892",X"F9C8",X"FB01",X"FC3E",X"FD7E",X"FEBE");

constant TblA : Tbl (0 to 255) := (X"0001",X"0001",X"1FFF",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001");

constant TblB : Tbl (0 to 255) := (X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"1FFF",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001");

constant TblC : Tbl (0 to 255) := (X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"1FFF",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001");

constant TblD : Tbl (0 to 255) := (X"1FFF",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001");

constant TblE : Tbl (0 to 255) := (X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",
X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"1FFF",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001");

begin

    process(clk,raz)
    begin
        if(raz='0')then 
            i <= 0;
            Write <= (others => '1');
            Reuse <= (others => '0');
            ect <= e00;
            
        elsif(clk'event and clk='1')then

            case ect is

                when e00 =>
                    Write <= (others => '0');
                    ect <= e0;                                  

                when e0 =>                    
                    if(i=255)then
                        Write <= (others => '1');
                        Reuse <= (others => '1');
                        ect <= eX;
                    else
                        i <= i+1;
                        ect <= e0;
                    end if;

                when eX =>
                    null; 

            end case;
        end if;
    end process;

data <= TblE(i) & TblD(i) & TblC(i) & TblB(i) & TblA(i);

end architecture;