------------------------------------------------------------------------------
--  This file is a part of the LPP VHDL IP LIBRARY
--  Copyright (C) 2009 - 2010, Laboratory of Plasmas Physic - CNRS
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
-------------------------------------------------------------------------------
--                    Author : Alexis Jeandet
--                     Mail : alexis.jeandet@lpp.polytechnique.fr
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use std.textio.all;
  


package lpp_amba is

component APB_ADVANCED_TRIGGER is
  generic (
    pindex   : integer := 0;
    paddr    : integer := 0
    );
  port (
    rstn   : in  std_ulogic;
    clk    : in  std_ulogic;
    apbi   : in  apb_slv_in_type;
    apbo   : out apb_slv_out_type;
    
    SPW_Tickout : IN STD_LOGIC;
    CoarseTime  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    FineTime    : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

    Trigger     : OUT STD_LOGIC
    );
end component;

component APB_ADVANCED_TRIGGER_v is
  generic (
    pindex   : integer;
    paddr    : integer;
    count    : integer range 1 to 8 := 1
  );
  port (
    rstn   : in  std_ulogic;
    clk    : in  std_ulogic;
    apbi   : in  apb_slv_in_type;
    apbo   : out apb_slv_out_type;

    SPW_Tickout : IN STD_LOGIC;
    CoarseTime  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    FineTime    : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

    Trigger     : OUT STD_LOGIC_VECTOR(count-1 DOWNTO 0)
    );
end component;

component APB_SIMPLE_DIODE is
  generic (
    pindex   : integer := 0;
    paddr    : integer := 0;
    pmask    : integer := 16#fff#;
    pirq     : integer := 0;
    abits    : integer := 8);
  port (
    rst    : in  std_ulogic;
    clk    : in  std_ulogic;
    apbi   : in  apb_slv_in_type;
    apbo   : out apb_slv_out_type;
    LED    : out std_ulogic
    );
end component;


component APB_MULTI_DIODE is
  generic (
    pindex   : integer := 0;
    paddr    : integer := 0;
    pmask    : integer := 16#fff#;
    pirq     : integer := 0;
    abits    : integer := 8);
  port (
    rst    : in  std_ulogic;
    clk    : in  std_ulogic;
    apbi   : in  apb_slv_in_type;
    apbo   : out apb_slv_out_type;
    LED    : out std_logic_vector(2 downto 0)
    );
end component;

end;
