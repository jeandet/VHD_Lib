-- Version: 9.1 SP5 9.1.5.1

library ieee;
use ieee.std_logic_1164.all;
library Axcelerator;
use Axcelerator.all;

entity actar is 
    port( DataA : in std_logic_vector(15 downto 0); DataB : in 
        std_logic_vector(15 downto 0); Mult : out 
        std_logic_vector(31 downto 0);Clock : in std_logic) ;
end actar;


architecture DEF_ARCH of  actar is

    component DF1
        port(D, CLK : in std_logic := 'U'; Q : out std_logic) ;
    end component;

    component XOR2
        port(A, B : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AO6
        port(A, B, C, D : in std_logic := 'U'; Y : out std_logic
        ) ;
    end component;

    component FA1
        port(A, B, CI : in std_logic := 'U'; CO, S : out 
        std_logic) ;
    end component;

    component MX2
        port(A, B, S : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component ADD1
        port(A, B, FCI : in std_logic := 'U'; S, FCO : out 
        std_logic) ;
    end component;

    component BUFF
        port(A : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component HA1
        port(A, B : in std_logic := 'U'; CO, S : out std_logic) ;
    end component;

    component OR3
        port(A, B, C : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AND3
        port(A, B, C : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AO16
        port(A, B, C : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AO1
        port(A, B, C : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AND2
        port(A, B : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component FCINIT_BUFF
        port(A : in std_logic := 'U'; FCO : out std_logic) ;
    end component;

    component AND2A
        port(A, B : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component AOI1
        port(A, B, C : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    component FCEND_BUFF
        port(FCI : in std_logic := 'U'; CO : out std_logic) ;
    end component;

    component VCC
        port( Y : out std_logic);
    end component;

    component GND
        port( Y : out std_logic);
    end component;

    signal S_0_net, S_1_net, S_2_net, S_3_net, S_4_net, S_5_net, 
        S_6_net, S_7_net, E_0_net, E_1_net, E_2_net, E_3_net, 
        E_4_net, E_5_net, E_6_net, E_7_net, EBAR, PP0_0_net, 
        PP0_1_net, PP0_2_net, PP0_3_net, PP0_4_net, PP0_5_net, 
        PP0_6_net, PP0_7_net, PP0_8_net, PP0_9_net, PP0_10_net, 
        PP0_11_net, PP0_12_net, PP0_13_net, PP0_14_net, 
        PP0_15_net, PP0_16_net, PP1_0_net, PP1_1_net, PP1_2_net, 
        PP1_3_net, PP1_4_net, PP1_5_net, PP1_6_net, PP1_7_net, 
        PP1_8_net, PP1_9_net, PP1_10_net, PP1_11_net, PP1_12_net, 
        PP1_13_net, PP1_14_net, PP1_15_net, PP1_16_net, PP2_0_net, 
        PP2_1_net, PP2_2_net, PP2_3_net, PP2_4_net, PP2_5_net, 
        PP2_6_net, PP2_7_net, PP2_8_net, PP2_9_net, PP2_10_net, 
        PP2_11_net, PP2_12_net, PP2_13_net, PP2_14_net, 
        PP2_15_net, PP2_16_net, PP3_0_net, PP3_1_net, PP3_2_net, 
        PP3_3_net, PP3_4_net, PP3_5_net, PP3_6_net, PP3_7_net, 
        PP3_8_net, PP3_9_net, PP3_10_net, PP3_11_net, PP3_12_net, 
        PP3_13_net, PP3_14_net, PP3_15_net, PP3_16_net, PP4_0_net, 
        PP4_1_net, PP4_2_net, PP4_3_net, PP4_4_net, PP4_5_net, 
        PP4_6_net, PP4_7_net, PP4_8_net, PP4_9_net, PP4_10_net, 
        PP4_11_net, PP4_12_net, PP4_13_net, PP4_14_net, 
        PP4_15_net, PP4_16_net, PP5_0_net, PP5_1_net, PP5_2_net, 
        PP5_3_net, PP5_4_net, PP5_5_net, PP5_6_net, PP5_7_net, 
        PP5_8_net, PP5_9_net, PP5_10_net, PP5_11_net, PP5_12_net, 
        PP5_13_net, PP5_14_net, PP5_15_net, PP5_16_net, PP6_0_net, 
        PP6_1_net, PP6_2_net, PP6_3_net, PP6_4_net, PP6_5_net, 
        PP6_6_net, PP6_7_net, PP6_8_net, PP6_9_net, PP6_10_net, 
        PP6_11_net, PP6_12_net, PP6_13_net, PP6_14_net, 
        PP6_15_net, PP6_16_net, PP7_0_net, PP7_1_net, PP7_2_net, 
        PP7_3_net, PP7_4_net, PP7_5_net, PP7_6_net, PP7_7_net, 
        PP7_8_net, PP7_9_net, PP7_10_net, PP7_11_net, PP7_12_net, 
        PP7_13_net, PP7_14_net, PP7_15_net, PP7_16_net, 
        SumA_0_net, SumA_1_net, SumA_2_net, SumA_3_net, 
        SumA_4_net, SumA_5_net, SumA_6_net, SumA_7_net, 
        SumA_8_net, SumA_9_net, SumA_10_net, SumA_11_net, 
        SumA_12_net, SumA_13_net, SumA_14_net, SumA_15_net, 
        SumA_16_net, SumA_17_net, SumA_18_net, SumA_19_net, 
        SumA_20_net, SumA_21_net, SumA_22_net, SumA_23_net, 
        SumA_24_net, SumA_25_net, SumA_26_net, SumA_27_net, 
        SumA_28_net, SumA_29_net, SumA_30_net, SumB_0_net, 
        SumB_1_net, SumB_2_net, SumB_3_net, SumB_4_net, 
        SumB_5_net, SumB_6_net, SumB_7_net, SumB_8_net, 
        SumB_9_net, SumB_10_net, SumB_11_net, SumB_12_net, 
        SumB_13_net, SumB_14_net, SumB_15_net, SumB_16_net, 
        SumB_17_net, SumB_18_net, SumB_19_net, SumB_20_net, 
        SumB_21_net, SumB_22_net, SumB_23_net, SumB_24_net, 
        SumB_25_net, SumB_26_net, SumB_27_net, SumB_28_net, 
        SumB_29_net, SumB_30_net, DF1_117_Q, DF1_114_Q, DF1_25_Q, 
        DF1_111_Q, DF1_143_Q, DF1_124_Q, DF1_18_Q, DF1_30_Q, 
        DF1_97_Q, DF1_90_Q, DF1_102_Q, DF1_63_Q, DF1_140_Q, 
        DF1_137_Q, DF1_45_Q, DF1_73_Q, DF1_23_Q, DF1_120_Q, 
        DF1_36_Q, DF1_130_Q, DF1_42_Q, DF1_8_Q, DF1_79_Q, 
        DF1_78_Q, DF1_135_Q, DF1_20_Q, DF1_112_Q, DF1_61_Q, 
        DF1_123_Q, DF1_70_Q, DF1_55_Q, DF1_28_Q, DF1_95_Q, 
        DF1_94_Q, DF1_2_Q, DF1_34_Q, DF1_125_Q, DF1_77_Q, 
        DF1_145_Q, DF1_88_Q, DF1_49_Q, DF1_17_Q, DF1_85_Q, 
        DF1_84_Q, DF1_147_Q, DF1_27_Q, DF1_115_Q, DF1_66_Q, 
        DF1_133_Q, DF1_76_Q, DF1_10_Q, DF1_127_Q, DF1_51_Q, 
        DF1_50_Q, DF1_107_Q, DF1_144_Q, DF1_81_Q, DF1_33_Q, 
        DF1_98_Q, DF1_43_Q, DF1_122_Q, DF1_96_Q, DF1_13_Q, 
        DF1_11_Q, DF1_67_Q, DF1_106_Q, DF1_48_Q, DF1_151_Q, 
        DF1_58_Q, DF1_6_Q, DF1_103_Q, DF1_64_Q, DF1_141_Q, 
        DF1_138_Q, DF1_46_Q, DF1_74_Q, DF1_24_Q, DF1_121_Q, 
        DF1_37_Q, DF1_131_Q, DF1_59_Q, DF1_31_Q, DF1_100_Q, 
        DF1_99_Q, DF1_5_Q, DF1_41_Q, DF1_132_Q, DF1_82_Q, 
        DF1_150_Q, DF1_91_Q, DF1_101_Q, DF1_62_Q, DF1_139_Q, 
        DF1_136_Q, DF1_44_Q, DF1_72_Q, DF1_22_Q, DF1_119_Q, 
        DF1_35_Q, DF1_129_Q, DF1_68_Q, DF1_118_Q, DF1_16_Q, 
        DF1_3_Q, DF1_86_Q, DF1_109_Q, DF1_60_Q, DF1_83_Q, 
        DF1_54_Q, DF1_53_Q, DF1_19_Q, DF1_69_Q, DF1_113_Q, 
        DF1_105_Q, DF1_38_Q, DF1_56_Q, DF1_12_Q, DF1_32_Q, 
        DF1_4_Q, DF1_1_Q, DF1_152_Q, DF1_52_Q, DF1_93_Q, DF1_80_Q, 
        DF1_14_Q, DF1_39_Q, DF1_146_Q, DF1_9_Q, DF1_134_Q, 
        DF1_126_Q, DF1_7_Q, DF1_57_Q, DF1_104_Q, DF1_89_Q, 
        DF1_26_Q, DF1_47_Q, DF1_0_Q, DF1_21_Q, DF1_148_Q, 
        DF1_142_Q, DF1_92_Q, DF1_149_Q, DF1_40_Q, DF1_29_Q, 
        DF1_110_Q, DF1_128_Q, DF1_87_Q, DF1_108_Q, DF1_75_Q, 
        DF1_71_Q, DF1_65_Q, DF1_116_Q, DF1_15_Q, HA1_13_S, 
        HA1_13_CO, FA1_94_S, FA1_94_CO, FA1_63_S, FA1_63_CO, 
        HA1_0_S, HA1_0_CO, FA1_71_S, FA1_71_CO, FA1_26_S, 
        FA1_26_CO, FA1_42_S, FA1_42_CO, FA1_24_S, FA1_24_CO, 
        HA1_12_S, HA1_12_CO, FA1_43_S, FA1_43_CO, FA1_90_S, 
        FA1_90_CO, HA1_6_S, HA1_6_CO, FA1_41_S, FA1_41_CO, 
        FA1_83_S, FA1_83_CO, HA1_9_S, HA1_9_CO, FA1_85_S, 
        FA1_85_CO, FA1_10_S, FA1_10_CO, HA1_2_S, HA1_2_CO, 
        FA1_67_S, FA1_67_CO, FA1_6_S, FA1_6_CO, HA1_1_S, HA1_1_CO, 
        FA1_86_S, FA1_86_CO, FA1_55_S, FA1_55_CO, FA1_3_S, 
        FA1_3_CO, HA1_8_S, HA1_8_CO, HA1_7_S, HA1_7_CO, FA1_30_S, 
        FA1_30_CO, FA1_29_S, FA1_29_CO, HA1_15_S, HA1_15_CO, 
        FA1_28_S, FA1_28_CO, FA1_14_S, FA1_14_CO, FA1_89_S, 
        FA1_89_CO, FA1_62_S, FA1_62_CO, FA1_5_S, FA1_5_CO, 
        FA1_12_S, FA1_12_CO, FA1_9_S, FA1_9_CO, FA1_38_S, 
        FA1_38_CO, FA1_37_S, FA1_37_CO, FA1_87_S, FA1_87_CO, 
        FA1_34_S, FA1_34_CO, FA1_44_S, FA1_44_CO, FA1_13_S, 
        FA1_13_CO, FA1_77_S, FA1_77_CO, FA1_33_S, FA1_33_CO, 
        FA1_40_S, FA1_40_CO, FA1_36_S, FA1_36_CO, FA1_61_S, 
        FA1_61_CO, FA1_60_S, FA1_60_CO, FA1_11_S, FA1_11_CO, 
        FA1_56_S, FA1_56_CO, FA1_27_S, FA1_27_CO, FA1_1_S, 
        FA1_1_CO, FA1_68_S, FA1_68_CO, FA1_18_S, FA1_18_CO, 
        FA1_22_S, FA1_22_CO, FA1_21_S, FA1_21_CO, FA1_51_S, 
        FA1_51_CO, FA1_50_S, FA1_50_CO, HA1_14_S, HA1_14_CO, 
        FA1_47_S, FA1_47_CO, HA1_10_S, HA1_10_CO, HA1_11_S, 
        HA1_11_CO, FA1_75_S, FA1_75_CO, FA1_31_S, FA1_31_CO, 
        FA1_35_S, FA1_35_CO, FA1_32_S, FA1_32_CO, FA1_58_S, 
        FA1_58_CO, FA1_57_S, FA1_57_CO, FA1_7_S, FA1_7_CO, 
        FA1_54_S, FA1_54_CO, FA1_25_S, FA1_25_CO, FA1_0_S, 
        FA1_0_CO, FA1_66_S, FA1_66_CO, FA1_15_S, FA1_15_CO, 
        FA1_20_S, FA1_20_CO, FA1_17_S, FA1_17_CO, FA1_49_S, 
        FA1_49_CO, FA1_48_S, FA1_48_CO, FA1_92_S, FA1_92_CO, 
        FA1_45_S, FA1_45_CO, FA1_70_S, FA1_70_CO, FA1_52_S, 
        FA1_52_CO, FA1_8_S, FA1_8_CO, FA1_65_S, FA1_65_CO, 
        HA1_5_S, HA1_5_CO, FA1_74_CO, FA1_74_S, HA1_3_CO, HA1_3_S, 
        FA1_78_CO, FA1_78_S, FA1_72_CO, FA1_72_S, HA1_4_CO, 
        HA1_4_S, FA1_73_CO, FA1_73_S, FA1_39_CO, FA1_39_S, 
        FA1_81_CO, FA1_81_S, FA1_2_CO, FA1_2_S, FA1_16_CO, 
        FA1_16_S, FA1_91_CO, FA1_91_S, FA1_93_CO, FA1_93_S, 
        FA1_88_CO, FA1_88_S, FA1_76_CO, FA1_76_S, FA1_82_CO, 
        FA1_82_S, FA1_95_CO, FA1_95_S, FA1_84_CO, FA1_84_S, 
        FA1_4_CO, FA1_4_S, FA1_46_CO, FA1_46_S, FA1_96_CO, 
        FA1_96_S, FA1_59_CO, FA1_59_S, FA1_80_CO, FA1_80_S, 
        FA1_69_CO, FA1_69_S, FA1_53_CO, FA1_53_S, FA1_79_CO, 
        FA1_79_S, FA1_64_CO, FA1_64_S, FA1_23_CO, FA1_23_S, 
        FA1_19_CO, FA1_19_S, BUF_29_Y, BUF_8_Y, BUF_21_Y, 
        BUF_35_Y, BUF_27_Y, BUF_25_Y, BUF_28_Y, BUF_4_Y, BUF_39_Y, 
        BUF_2_Y, BUF_45_Y, BUF_36_Y, BUF_7_Y, BUF_13_Y, BUF_5_Y, 
        BUF_44_Y, BUF_14_Y, BUF_19_Y, BUF_10_Y, BUF_38_Y, 
        BUF_43_Y, BUF_9_Y, BUF_42_Y, BUF_15_Y, BUF_24_Y, BUF_1_Y, 
        BUF_16_Y, BUF_32_Y, BUF_0_Y, BUF_31_Y, BUF_46_Y, BUF_40_Y, 
        BUF_47_Y, BUF_41_Y, XOR2_24_Y, XOR2_19_Y, AO1_4_Y, 
        XOR2_6_Y, AO16_2_Y, AO6_57_Y, AO6_107_Y, AO6_104_Y, 
        AO6_82_Y, MX2_3_Y, AO6_115_Y, AO6_13_Y, AO6_42_Y, 
        XOR2_29_Y, AO16_4_Y, AO6_25_Y, AO6_36_Y, AO6_65_Y, 
        AND2_6_Y, AO6_28_Y, AO6_50_Y, AO6_72_Y, AO6_60_Y, 
        AO6_52_Y, OR3_3_Y, AND3_5_Y, BUF_17_Y, BUF_6_Y, XOR2_1_Y, 
        XOR2_7_Y, AO1_6_Y, XOR2_3_Y, AO16_8_Y, AO6_91_Y, AO6_93_Y, 
        AO6_56_Y, AO6_54_Y, MX2_5_Y, AO6_74_Y, AO6_102_Y, AO6_3_Y, 
        XOR2_8_Y, AO16_5_Y, AO6_44_Y, AO6_0_Y, AO6_97_Y, AND2_3_Y, 
        AO6_40_Y, AO6_67_Y, AO6_64_Y, AO6_90_Y, AO6_55_Y, OR3_0_Y, 
        AND3_3_Y, BUF_18_Y, BUF_11_Y, XOR2_27_Y, XOR2_13_Y, 
        AO1_5_Y, XOR2_4_Y, AO16_3_Y, AO6_23_Y, AO6_113_Y, 
        AO6_22_Y, AO6_1_Y, MX2_1_Y, AO6_78_Y, AO6_84_Y, AO6_33_Y, 
        XOR2_25_Y, AO16_13_Y, AO6_105_Y, AO6_46_Y, AO6_61_Y, 
        AND2_2_Y, AO6_68_Y, AO6_35_Y, AO6_29_Y, AO6_98_Y, 
        AO6_66_Y, OR3_2_Y, AND3_6_Y, BUF_26_Y, BUF_23_Y, 
        XOR2_16_Y, XOR2_26_Y, AND2A_1_Y, AO6_88_Y, AO6_51_Y, 
        AO6_48_Y, AO6_41_Y, MX2_2_Y, AO6_30_Y, AO6_92_Y, AO6_11_Y, 
        AND2A_0_Y, AO6_76_Y, AO6_73_Y, AO6_114_Y, AND2_0_Y, 
        AO6_63_Y, AO6_32_Y, AO6_45_Y, AO6_38_Y, AO6_4_Y, OR3_1_Y, 
        AND3_1_Y, BUF_22_Y, BUF_20_Y, XOR2_12_Y, XOR2_11_Y, 
        AO1_3_Y, XOR2_18_Y, AO16_6_Y, AO6_69_Y, AO6_21_Y, 
        AO6_34_Y, AO6_6_Y, MX2_4_Y, AO6_95_Y, AO6_101_Y, 
        AO6_117_Y, XOR2_2_Y, AO16_12_Y, AO6_109_Y, AO6_7_Y, 
        AO6_14_Y, AND2_7_Y, AO6_31_Y, AO6_111_Y, AO6_118_Y, 
        AO6_2_Y, AO6_96_Y, OR3_4_Y, AND3_7_Y, BUF_37_Y, BUF_33_Y, 
        XOR2_0_Y, XOR2_20_Y, AO1_0_Y, XOR2_5_Y, AO16_0_Y, 
        AO6_75_Y, AO6_53_Y, AO6_20_Y, AO6_49_Y, MX2_6_Y, AO6_94_Y, 
        AO6_87_Y, AO6_37_Y, XOR2_10_Y, AO16_1_Y, AO6_89_Y, 
        AO6_83_Y, AO6_10_Y, AND2_4_Y, AO6_85_Y, AO6_71_Y, 
        AO6_58_Y, AO6_26_Y, AO6_112_Y, OR3_7_Y, AND3_0_Y, 
        BUF_12_Y, BUF_3_Y, XOR2_14_Y, XOR2_15_Y, AO1_1_Y, 
        XOR2_28_Y, AO16_7_Y, AO6_15_Y, AO6_59_Y, AO6_12_Y, 
        AO6_86_Y, MX2_7_Y, AO6_8_Y, AO6_99_Y, AO6_100_Y, 
        XOR2_17_Y, AO16_11_Y, AO6_103_Y, AO6_43_Y, AO6_16_Y, 
        AND2_5_Y, AO6_110_Y, AO6_62_Y, AO6_108_Y, AO6_70_Y, 
        AO6_18_Y, OR3_5_Y, AND3_4_Y, BUF_34_Y, BUF_30_Y, XOR2_9_Y, 
        XOR2_22_Y, AO1_2_Y, XOR2_23_Y, AO16_9_Y, AO6_79_Y, 
        AO6_5_Y, AO6_119_Y, AO6_116_Y, MX2_0_Y, AO6_39_Y, 
        AO6_81_Y, AO6_17_Y, XOR2_21_Y, AO16_10_Y, AO6_9_Y, 
        AO6_77_Y, AO6_24_Y, AND2_1_Y, AO6_80_Y, AO6_27_Y, 
        AO6_106_Y, AO6_47_Y, AO6_19_Y, OR3_6_Y, AND3_2_Y, 
        FCEND_BUFF_0_CO, FCINIT_BUFF_0_FCO, ADD1_Mult_1_FCO, 
        ADD1_Mult_2_FCO, ADD1_Mult_3_FCO, ADD1_Mult_4_FCO, 
        ADD1_Mult_5_FCO, ADD1_Mult_6_FCO, ADD1_Mult_7_FCO, 
        ADD1_Mult_8_FCO, ADD1_Mult_9_FCO, ADD1_Mult_10_FCO, 
        ADD1_Mult_11_FCO, ADD1_Mult_12_FCO, ADD1_Mult_13_FCO, 
        ADD1_Mult_14_FCO, ADD1_Mult_15_FCO, ADD1_Mult_16_FCO, 
        ADD1_Mult_17_FCO, ADD1_Mult_18_FCO, ADD1_Mult_19_FCO, 
        ADD1_Mult_20_FCO, ADD1_Mult_21_FCO, ADD1_Mult_22_FCO, 
        ADD1_Mult_23_FCO, ADD1_Mult_24_FCO, ADD1_Mult_25_FCO, 
        ADD1_Mult_26_FCO, ADD1_Mult_27_FCO, ADD1_Mult_28_FCO, 
        ADD1_Mult_29_FCO, ADD1_Mult_30_FCO, ADD1_Mult_31_FCO, 
        VCC_1_net, GND_1_net : std_logic ;
    begin   

    VCC_2_net : VCC port map(Y => VCC_1_net);
    GND_2_net : GND port map(Y => GND_1_net);
    DF1_SumB_0_inst : DF1
      port map(D => DF1_0_Q, CLK => Clock, Q => SumB_0_net);
    XOR2_PP7_9_inst : XOR2
      port map(A => AO6_6_Y, B => BUF_20_Y, Y => PP7_9_net);
    DF1_145 : DF1
      port map(D => PP2_4_net, CLK => Clock, Q => DF1_145_Q);
    DF1_SumA_17_inst : DF1
      port map(D => FA1_93_CO, CLK => Clock, Q => SumA_17_net);
    AO6_7 : AO6
      port map(A => BUF_4_Y, B => AO16_12_Y, C => BUF_2_Y, D => 
        XOR2_2_Y, Y => AO6_7_Y);
    DF1_60 : DF1
      port map(D => PP6_4_net, CLK => Clock, Q => DF1_60_Q);
    FA1_33 : FA1
      port map(A => FA1_90_CO, B => HA1_6_CO, CI => FA1_83_S, 
        CO => FA1_33_CO, S => FA1_33_S);
    FA1_46 : FA1
      port map(A => HA1_11_CO, B => DF1_127_Q, CI => FA1_75_S, 
        CO => FA1_46_CO, S => FA1_46_S);
    DF1_SumA_6_inst : DF1
      port map(D => FA1_46_CO, CLK => Clock, Q => SumA_6_net);
    MX2_PP1_16_inst : MX2
      port map(A => MX2_1_Y, B => AO1_5_Y, S => AO16_3_Y, Y => 
        PP1_16_net);
    DF1_65 : DF1
      port map(D => E_6_net, CLK => Clock, Q => DF1_65_Q);
    ADD1_Mult_23_inst : ADD1
      port map(A => SumA_22_net, B => SumB_22_net, FCI => 
        ADD1_Mult_22_FCO, S => Mult(23), FCO => ADD1_Mult_23_FCO);
    DF1_SumB_6_inst : DF1
      port map(D => FA1_81_S, CLK => Clock, Q => SumB_6_net);
    FA1_86 : FA1
      port map(A => DF1_106_Q, B => VCC_1_net, CI => DF1_72_Q, 
        CO => FA1_86_CO, S => FA1_86_S);
    DF1_SumB_13_inst : DF1
      port map(D => FA1_96_S, CLK => Clock, Q => SumB_13_net);
    FA1_44 : FA1
      port map(A => FA1_71_CO, B => HA1_12_S, CI => FA1_42_S, 
        CO => FA1_44_CO, S => FA1_44_S);
    FA1_9 : FA1
      port map(A => DF1_40_Q, B => DF1_150_Q, CI => FA1_94_CO, 
        CO => FA1_9_CO, S => FA1_9_S);
    FA1_90 : FA1
      port map(A => DF1_96_Q, B => DF1_28_Q, CI => DF1_62_Q, 
        CO => FA1_90_CO, S => FA1_90_S);
    DF1_SumA_22_inst : DF1
      port map(D => FA1_74_CO, CLK => Clock, Q => SumA_22_net);
    BUF_36 : BUFF
      port map(A => DataA(5), Y => BUF_36_Y);
    AO6_30 : AO6
      port map(A => BUF_16_Y, B => AND2A_1_Y, C => BUF_0_Y, D => 
        DataB(0), Y => AO6_30_Y);
    DF1_SumB_4_inst : DF1
      port map(D => FA1_82_S, CLK => Clock, Q => SumB_4_net);
    XOR2_PP0_13_inst : XOR2
      port map(A => AO6_51_Y, B => BUF_23_Y, Y => PP0_13_net);
    XOR2_PP5_4_inst : XOR2
      port map(A => AO6_36_Y, B => BUF_47_Y, Y => PP5_4_net);
    AO6_8 : AO6
      port map(A => BUF_16_Y, B => AO16_7_Y, C => BUF_0_Y, D => 
        XOR2_28_Y, Y => AO6_8_Y);
    FA1_84 : FA1
      port map(A => DF1_130_Q, B => DF1_143_Q, CI => DF1_2_Q, 
        CO => FA1_84_CO, S => FA1_84_S);
    HA1_11 : HA1
      port map(A => DF1_42_Q, B => DF1_124_Q, CO => HA1_11_CO, 
        S => HA1_11_S);
    XOR2_PP6_6_inst : XOR2
      port map(A => AO6_44_Y, B => BUF_17_Y, Y => PP6_6_net);
    AO6_25 : AO6
      port map(A => BUF_36_Y, B => AO16_4_Y, C => BUF_13_Y, D => 
        XOR2_29_Y, Y => AO6_25_Y);
    FA1_63 : FA1
      port map(A => DF1_123_Q, B => DF1_137_Q, CI => DF1_84_Q, 
        CO => FA1_63_CO, S => FA1_63_S);
    AO6_51 : AO6
      port map(A => BUF_24_Y, B => AND2A_1_Y, C => BUF_16_Y, D => 
        DataB(0), Y => AO6_51_Y);
    FA1_75 : FA1
      port map(A => DF1_8_Q, B => DF1_18_Q, CI => DF1_125_Q, 
        CO => FA1_75_CO, S => FA1_75_S);
    AO6_16 : AO6
      port map(A => BUF_29_Y, B => AO16_11_Y, C => BUF_21_Y, D => 
        XOR2_17_Y, Y => AO6_16_Y);
    XOR2_PP6_4_inst : XOR2
      port map(A => AO6_0_Y, B => BUF_17_Y, Y => PP6_4_net);
    XOR2_PP6_10_inst : XOR2
      port map(A => AO6_56_Y, B => BUF_6_Y, Y => PP6_10_net);
    XOR2_PP5_13_inst : XOR2
      port map(A => AO6_107_Y, B => BUF_41_Y, Y => PP5_13_net);
    DF1_SumA_30_inst : DF1
      port map(D => DF1_116_Q, CLK => Clock, Q => SumA_30_net);
    DF1_88 : DF1
      port map(D => PP2_5_net, CLK => Clock, Q => DF1_88_Q);
    OR3_6 : OR3
      port map(A => DataB(3), B => DataB(4), C => DataB(5), Y => 
        OR3_6_Y);
    DF1_SumB_5_inst : DF1
      port map(D => FA1_46_S, CLK => Clock, Q => SumB_5_net);
    FA1_26 : FA1
      port map(A => DF1_43_Q, B => DF1_70_Q, CI => DF1_91_Q, 
        CO => FA1_26_CO, S => FA1_26_S);
    BUF_43 : BUFF
      port map(A => DataA(10), Y => BUF_43_Y);
    DF1_134 : DF1
      port map(D => PP7_9_net, CLK => Clock, Q => DF1_134_Q);
    DF1_13 : DF1
      port map(D => PP3_11_net, CLK => Clock, Q => DF1_13_Q);
    ADD1_Mult_28_inst : ADD1
      port map(A => SumA_27_net, B => SumB_27_net, FCI => 
        ADD1_Mult_27_FCO, S => Mult(28), FCO => ADD1_Mult_28_FCO);
    XOR2_PP2_4_inst : XOR2
      port map(A => AO6_77_Y, B => BUF_34_Y, Y => PP2_4_net);
    FA1_24 : FA1
      port map(A => DF1_122_Q, B => DF1_55_Q, CI => DF1_101_Q, 
        CO => FA1_24_CO, S => FA1_24_S);
    MX2_1 : MX2
      port map(A => BUF_11_Y, B => XOR2_13_Y, S => XOR2_4_Y, Y => 
        MX2_1_Y);
    ADD1_Mult_6_inst : ADD1
      port map(A => SumA_5_net, B => SumB_5_net, FCI => 
        ADD1_Mult_5_FCO, S => Mult(6), FCO => ADD1_Mult_6_FCO);
    AO6_35 : AO6
      port map(A => BUF_39_Y, B => AO16_13_Y, C => BUF_45_Y, D => 
        XOR2_25_Y, Y => AO6_35_Y);
    AO6_74 : AO6
      port map(A => BUF_32_Y, B => AO16_8_Y, C => BUF_31_Y, D => 
        XOR2_3_Y, Y => AO6_74_Y);
    DF1_104 : DF1
      port map(D => PP7_13_net, CLK => Clock, Q => DF1_104_Q);
    XOR2_PP2_11_inst : XOR2
      port map(A => AO6_81_Y, B => BUF_30_Y, Y => PP2_11_net);
    DF1_10 : DF1
      port map(D => PP2_16_net, CLK => Clock, Q => DF1_10_Q);
    DF1_33 : DF1
      port map(D => PP3_6_net, CLK => Clock, Q => DF1_33_Q);
    AO6_108 : AO6
      port map(A => BUF_21_Y, B => AO16_11_Y, C => BUF_27_Y, D => 
        XOR2_17_Y, Y => AO6_108_Y);
    FA1_51 : FA1
      port map(A => DF1_105_Q, B => DF1_99_Q, CI => HA1_8_CO, 
        CO => FA1_51_CO, S => FA1_51_S);
    XOR2_PP1_15_inst : XOR2
      port map(A => AO6_23_Y, B => BUF_11_Y, Y => PP1_15_net);
    DF1_0 : DF1
      port map(D => S_0_net, CLK => Clock, Q => DF1_0_Q);
    DF1_9 : DF1
      port map(D => PP7_8_net, CLK => Clock, Q => DF1_9_Q);
    AO6_67 : AO6
      port map(A => BUF_2_Y, B => AO16_5_Y, C => BUF_36_Y, D => 
        XOR2_8_Y, Y => AO6_67_Y);
    BUF_15 : BUFF
      port map(A => DataA(11), Y => BUF_15_Y);
    AO6_2 : AO6
      port map(A => BUF_44_Y, B => AO16_12_Y, C => BUF_19_Y, D => 
        XOR2_2_Y, Y => AO6_2_Y);
    DF1_15 : DF1
      port map(D => EBAR, CLK => Clock, Q => DF1_15_Q);
    DF1_72 : DF1
      port map(D => PP5_10_net, CLK => Clock, Q => DF1_72_Q);
    DF1_41 : DF1
      port map(D => PP5_0_net, CLK => Clock, Q => DF1_41_Q);
    FA1_57 : FA1
      port map(A => FA1_28_CO, B => FA1_14_CO, CI => FA1_62_S, 
        CO => FA1_57_CO, S => FA1_57_S);
    BUF_25 : BUFF
      port map(A => DataA(2), Y => BUF_25_Y);
    DF1_30 : DF1
      port map(D => PP0_7_net, CLK => Clock, Q => DF1_30_Q);
    XOR2_PP4_7_inst : XOR2
      port map(A => AO6_85_Y, B => BUF_37_Y, Y => PP4_7_net);
    AO6_84 : AO6
      port map(A => BUF_43_Y, B => AO16_3_Y, C => BUF_42_Y, D => 
        XOR2_4_Y, Y => AO6_84_Y);
    FA1_0 : FA1
      port map(A => FA1_37_CO, B => FA1_87_CO, CI => FA1_44_S, 
        CO => FA1_0_CO, S => FA1_0_S);
    DF1_47 : DF1
      port map(D => PP7_16_net, CLK => Clock, Q => DF1_47_Q);
    FA1_15 : FA1
      port map(A => FA1_13_CO, B => FA1_77_CO, CI => FA1_40_S, 
        CO => FA1_15_CO, S => FA1_15_S);
    FA1_36 : FA1
      port map(A => FA1_83_CO, B => HA1_9_CO, CI => FA1_10_S, 
        CO => FA1_36_CO, S => FA1_36_S);
    XOR2_24 : XOR2
      port map(A => AND2_6_Y, B => BUF_47_Y, Y => XOR2_24_Y);
    DF1_35 : DF1
      port map(D => PP5_13_net, CLK => Clock, Q => DF1_35_Q);
    AO6_68 : AO6
      port map(A => BUF_7_Y, B => AO16_13_Y, C => BUF_5_Y, D => 
        XOR2_25_Y, Y => AO6_68_Y);
    XOR2_PP2_14_inst : XOR2
      port map(A => AO6_39_Y, B => BUF_30_Y, Y => PP2_14_net);
    FA1_34 : FA1
      port map(A => FA1_26_CO, B => DF1_29_Q, CI => FA1_24_S, 
        CO => FA1_34_CO, S => FA1_34_S);
    AO6_79 : AO6
      port map(A => BUF_0_Y, B => AO16_9_Y, C => BUF_46_Y, D => 
        XOR2_23_Y, Y => AO6_79_Y);
    BUF_16 : BUFF
      port map(A => DataA(13), Y => BUF_16_Y);
    DF1_SumA_7_inst : DF1
      port map(D => FA1_81_CO, CLK => Clock, Q => SumA_7_net);
    OR3_4 : OR3
      port map(A => DataB(13), B => DataB(14), C => DataB(15), 
        Y => OR3_4_Y);
    MX2_0 : MX2
      port map(A => BUF_30_Y, B => XOR2_22_Y, S => XOR2_23_Y, 
        Y => MX2_0_Y);
    AO6_3 : AO6
      port map(A => BUF_15_Y, B => AO16_8_Y, C => BUF_1_Y, D => 
        XOR2_3_Y, Y => AO6_3_Y);
    BUF_26 : BUFF
      port map(A => DataB(1), Y => BUF_26_Y);
    DF1_SumA_20_inst : DF1
      port map(D => FA1_2_CO, CLK => Clock, Q => SumA_20_net);
    AO6_115 : AO6
      port map(A => BUF_32_Y, B => AO16_2_Y, C => BUF_31_Y, D => 
        XOR2_6_Y, Y => AO6_115_Y);
    FA1_66 : FA1
      port map(A => FA1_34_CO, B => FA1_44_CO, CI => FA1_77_S, 
        CO => FA1_66_CO, S => FA1_66_S);
    FA1_45 : FA1
      port map(A => FA1_18_CO, B => FA1_22_CO, CI => FA1_51_S, 
        CO => FA1_45_CO, S => FA1_45_S);
    AO6_103 : AO6
      port map(A => BUF_45_Y, B => AO16_11_Y, C => BUF_7_Y, D => 
        XOR2_17_Y, Y => AO6_103_Y);
    AO6_89 : AO6
      port map(A => BUF_36_Y, B => AO16_1_Y, C => BUF_13_Y, D => 
        XOR2_10_Y, Y => AO6_89_Y);
    DF1_SumB_27_inst : DF1
      port map(D => FA1_19_S, CLK => Clock, Q => SumB_27_net);
    DF1_53 : DF1
      port map(D => PP6_7_net, CLK => Clock, Q => DF1_53_Q);
    HA1_8 : HA1
      port map(A => DF1_151_Q, B => VCC_1_net, CO => HA1_8_CO, 
        S => HA1_8_S);
    DF1_SumA_25_inst : DF1
      port map(D => FA1_69_CO, CLK => Clock, Q => SumA_25_net);
    FA1_85 : FA1
      port map(A => DF1_133_Q, B => DF1_15_Q, CI => DF1_37_Q, 
        CO => FA1_85_CO, S => FA1_85_S);
    FA1_64 : FA1
      port map(A => FA1_35_CO, B => FA1_29_S, CI => FA1_32_S, 
        CO => FA1_64_CO, S => FA1_64_S);
    XOR2_PP7_11_inst : XOR2
      port map(A => AO6_101_Y, B => BUF_20_Y, Y => PP7_11_net);
    XOR2_PP5_1_inst : XOR2
      port map(A => AO6_65_Y, B => BUF_47_Y, Y => PP5_1_net);
    DF1_50 : DF1
      port map(D => PP3_2_net, CLK => Clock, Q => DF1_50_Q);
    XOR2_PP4_10_inst : XOR2
      port map(A => AO6_20_Y, B => BUF_33_Y, Y => PP4_10_net);
    AO6_24 : AO6
      port map(A => BUF_29_Y, B => AO16_10_Y, C => BUF_21_Y, D => 
        XOR2_21_Y, Y => AO6_24_Y);
    XOR2_PP3_11_inst : XOR2
      port map(A => AO6_99_Y, B => BUF_3_Y, Y => PP3_11_net);
    XOR2_9 : XOR2
      port map(A => AND2_1_Y, B => BUF_34_Y, Y => XOR2_9_Y);
    XOR2_25 : XOR2
      port map(A => DataB(1), B => DataB(2), Y => XOR2_25_Y);
    DF1_24 : DF1
      port map(D => PP4_8_net, CLK => Clock, Q => DF1_24_Q);
    DF1_55 : DF1
      port map(D => PP1_13_net, CLK => Clock, Q => DF1_55_Q);
    FA1_7 : FA1
      port map(A => FA1_89_CO, B => FA1_62_CO, CI => FA1_12_S, 
        CO => FA1_7_CO, S => FA1_7_S);
    AND3_0 : AND3
      port map(A => DataB(7), B => DataB(8), C => DataB(9), Y => 
        AND3_0_Y);
    FA1_70 : FA1
      port map(A => FA1_51_CO, B => HA1_14_S, CI => FA1_21_CO, 
        CO => FA1_70_CO, S => FA1_70_S);
    XOR2_PP1_1_inst : XOR2
      port map(A => AO6_61_Y, B => BUF_18_Y, Y => PP1_1_net);
    AO16_4 : AO16
      port map(A => DataB(9), B => DataB(10), C => BUF_47_Y, Y => 
        AO16_4_Y);
    DF1_49 : DF1
      port map(D => PP2_6_net, CLK => Clock, Q => DF1_49_Q);
    MX2_7 : MX2
      port map(A => BUF_3_Y, B => XOR2_15_Y, S => XOR2_28_Y, Y => 
        MX2_7_Y);
    DF1_SumB_16_inst : DF1
      port map(D => FA1_93_S, CLK => Clock, Q => SumB_16_net);
    HA1_13 : HA1
      port map(A => DF1_112_Q, B => DF1_63_Q, CO => HA1_13_CO, 
        S => HA1_13_S);
    FA1_25 : FA1
      port map(A => FA1_9_CO, B => FA1_38_CO, CI => FA1_87_S, 
        CO => FA1_25_CO, S => FA1_25_S);
    XOR2_PP7_14_inst : XOR2
      port map(A => AO6_95_Y, B => BUF_20_Y, Y => PP7_14_net);
    DF1_86 : DF1
      port map(D => PP6_2_net, CLK => Clock, Q => DF1_86_Q);
    AO1_3 : AO1
      port map(A => XOR2_11_Y, B => OR3_4_Y, C => AND3_7_Y, Y => 
        AO1_3_Y);
    AND3_7 : AND3
      port map(A => DataB(13), B => DataB(14), C => DataB(15), 
        Y => AND3_7_Y);
    DF1_126 : DF1
      port map(D => PP7_10_net, CLK => Clock, Q => DF1_126_Q);
    OR3_0 : OR3
      port map(A => DataB(11), B => DataB(12), C => DataB(13), 
        Y => OR3_0_Y);
    MX2_6 : MX2
      port map(A => BUF_33_Y, B => XOR2_20_Y, S => XOR2_5_Y, Y => 
        MX2_6_Y);
    AO6_34 : AO6
      port map(A => BUF_38_Y, B => AO16_6_Y, C => BUF_9_Y, D => 
        XOR2_18_Y, Y => AO6_34_Y);
    XOR2_PP3_14_inst : XOR2
      port map(A => AO6_8_Y, B => BUF_3_Y, Y => PP3_14_net);
    AO16_1 : AO16
      port map(A => DataB(7), B => DataB(8), C => BUF_37_Y, Y => 
        AO16_1_Y);
    ADD1_Mult_10_inst : ADD1
      port map(A => SumA_9_net, B => SumB_9_net, FCI => 
        ADD1_Mult_9_FCO, S => Mult(10), FCO => ADD1_Mult_10_FCO);
    AO6_29 : AO6
      port map(A => BUF_21_Y, B => AO16_13_Y, C => BUF_27_Y, D => 
        XOR2_25_Y, Y => AO6_29_Y);
    XOR2_PP0_12_inst : XOR2
      port map(A => AO6_11_Y, B => BUF_23_Y, Y => PP0_12_net);
    DF1_SumB_18_inst : DF1
      port map(D => FA1_79_S, CLK => Clock, Q => SumB_18_net);
    AO1_0 : AO1
      port map(A => XOR2_20_Y, B => OR3_7_Y, C => AND3_0_Y, Y => 
        AO1_0_Y);
    DF1_SumB_7_inst : DF1
      port map(D => FA1_80_S, CLK => Clock, Q => SumB_7_net);
    DF1_149 : DF1
      port map(D => S_5_net, CLK => Clock, Q => DF1_149_Q);
    DF1_SumB_8_inst : DF1
      port map(D => FA1_64_S, CLK => Clock, Q => SumB_8_net);
    ADD1_Mult_16_inst : ADD1
      port map(A => SumA_15_net, B => SumB_15_net, FCI => 
        ADD1_Mult_15_FCO, S => Mult(16), FCO => ADD1_Mult_16_FCO);
    AO16_7 : AO16
      port map(A => DataB(5), B => DataB(6), C => BUF_3_Y, Y => 
        AO16_7_Y);
    DF1_64 : DF1
      port map(D => PP4_3_net, CLK => Clock, Q => DF1_64_Q);
    XOR2_18 : XOR2
      port map(A => DataB(13), B => DataB(14), Y => XOR2_18_Y);
    XOR2_PP5_12_inst : XOR2
      port map(A => AO6_42_Y, B => BUF_41_Y, Y => PP5_12_net);
    DF1_117 : DF1
      port map(D => PP0_0_net, CLK => Clock, Q => DF1_117_Q);
    XOR2_20 : XOR2
      port map(A => BUF_40_Y, B => DataB(9), Y => XOR2_20_Y);
    DF1_SumA_12_inst : DF1
      port map(D => FA1_76_CO, CLK => Clock, Q => SumA_12_net);
    FA1_1 : FA1
      port map(A => DF1_146_Q, B => DF1_22_Q, CI => FA1_86_CO, 
        CO => FA1_1_CO, S => FA1_1_S);
    FA1_35 : FA1
      port map(A => DF1_58_Q, B => DF1_50_Q, CI => HA1_7_CO, 
        CO => FA1_35_CO, S => FA1_35_S);
    FA1_53 : FA1
      port map(A => FA1_49_CO, B => FA1_1_S, CI => FA1_48_S, 
        CO => FA1_53_CO, S => FA1_53_S);
    MX2_PP3_16_inst : MX2
      port map(A => MX2_7_Y, B => AO1_1_Y, S => AO16_7_Y, Y => 
        PP3_16_net);
    FA1_10 : FA1
      port map(A => DF1_11_Q, B => DF1_94_Q, CI => DF1_136_Q, 
        CO => FA1_10_CO, S => FA1_10_S);
    AO6_39 : AO6
      port map(A => BUF_16_Y, B => AO16_9_Y, C => BUF_0_Y, D => 
        XOR2_23_Y, Y => AO6_39_Y);
    ADD1_Mult_30_inst : ADD1
      port map(A => SumA_29_net, B => SumB_29_net, FCI => 
        ADD1_Mult_29_FCO, S => Mult(30), FCO => ADD1_Mult_30_FCO);
    AO6_76 : AO6
      port map(A => BUF_45_Y, B => AND2A_0_Y, C => BUF_7_Y, D => 
        DataB(0), Y => AO6_76_Y);
    BUF_44 : BUFF
      port map(A => DataA(7), Y => BUF_44_Y);
    HA1_S_6_inst : HA1
      port map(A => XOR2_1_Y, B => DataB(13), CO => S_6_net, S => 
        PP6_0_net);
    DF1_28 : DF1
      port map(D => PP1_14_net, CLK => Clock, Q => DF1_28_Q);
    DF1_93 : DF1
      port map(D => PP7_3_net, CLK => Clock, Q => DF1_93_Q);
    AND2_4 : AND2
      port map(A => XOR2_10_Y, B => BUF_8_Y, Y => AND2_4_Y);
    AO6_61 : AO6
      port map(A => BUF_29_Y, B => AO16_13_Y, C => BUF_21_Y, D => 
        XOR2_25_Y, Y => AO6_61_Y);
    DF1_131 : DF1
      port map(D => PP4_11_net, CLK => Clock, Q => DF1_131_Q);
    MX2_PP6_16_inst : MX2
      port map(A => MX2_5_Y, B => AO1_6_Y, S => AO16_8_Y, Y => 
        PP6_16_net);
    XOR2_PP7_8_inst : XOR2
      port map(A => AO6_2_Y, B => BUF_22_Y, Y => PP7_8_net);
    ADD1_Mult_13_inst : ADD1
      port map(A => SumA_12_net, B => SumB_12_net, FCI => 
        ADD1_Mult_12_FCO, S => Mult(13), FCO => ADD1_Mult_13_FCO);
    AND2_0 : AND2
      port map(A => DataB(0), B => BUF_29_Y, Y => AND2_0_Y);
    DF1_90 : DF1
      port map(D => PP0_9_net, CLK => Clock, Q => DF1_90_Q);
    AO6_86 : AO6
      port map(A => BUF_14_Y, B => AO16_7_Y, C => BUF_10_Y, D => 
        XOR2_28_Y, Y => AO6_86_Y);
    DF1_110 : DF1
      port map(D => E_0_net, CLK => Clock, Q => DF1_110_Q);
    FA1_65 : FA1
      port map(A => DF1_32_Q, B => DF1_71_Q, CI => DF1_104_Q, 
        CO => FA1_65_CO, S => FA1_65_S);
    BUF_38 : BUFF
      port map(A => DataA(9), Y => BUF_38_Y);
    FA1_4 : FA1
      port map(A => FA1_15_CO, B => FA1_36_S, CI => FA1_20_S, 
        CO => FA1_4_CO, S => FA1_4_S);
    AO6_90 : AO6
      port map(A => BUF_44_Y, B => AO16_5_Y, C => BUF_19_Y, D => 
        XOR2_8_Y, Y => AO6_90_Y);
    AND2_6 : AND2
      port map(A => XOR2_29_Y, B => BUF_8_Y, Y => AND2_6_Y);
    XOR2_PP6_13_inst : XOR2
      port map(A => AO6_93_Y, B => BUF_6_Y, Y => PP6_13_net);
    DF1_101 : DF1
      port map(D => PP5_5_net, CLK => Clock, Q => DF1_101_Q);
    FA1_40 : FA1
      port map(A => FA1_43_CO, B => HA1_9_S, CI => FA1_41_S, 
        CO => FA1_40_CO, S => FA1_40_S);
    AO6_102 : AO6
      port map(A => BUF_9_Y, B => AO16_8_Y, C => BUF_15_Y, D => 
        XOR2_3_Y, Y => AO6_102_Y);
    DF1_95 : DF1
      port map(D => PP1_15_net, CLK => Clock, Q => DF1_95_Q);
    DF1_138 : DF1
      port map(D => PP4_5_net, CLK => Clock, Q => DF1_138_Q);
    DF1_SumA_29_inst : DF1
      port map(D => HA1_4_S, CLK => Clock, Q => SumA_29_net);
    AO6_107 : AO6
      port map(A => BUF_1_Y, B => AO16_2_Y, C => BUF_32_Y, D => 
        XOR2_6_Y, Y => AO6_107_Y);
    FA1_8 : FA1
      port map(A => DF1_57_Q, B => DF1_12_Q, CI => HA1_10_S, 
        CO => FA1_8_CO, S => FA1_8_S);
    FA1_80 : FA1
      port map(A => FA1_31_CO, B => FA1_30_S, CI => FA1_35_S, 
        CO => FA1_80_CO, S => FA1_80_S);
    DF1_81 : DF1
      port map(D => PP3_5_net, CLK => Clock, Q => DF1_81_Q);
    DF1_151 : DF1
      port map(D => PP3_16_net, CLK => Clock, Q => DF1_151_Q);
    XOR2_PP0_5_inst : XOR2
      port map(A => AO6_32_Y, B => BUF_26_Y, Y => PP0_5_net);
    HA1_5 : HA1
      port map(A => DF1_4_Q, B => VCC_1_net, CO => HA1_5_CO, S => 
        HA1_5_S);
    DF1_7 : DF1
      port map(D => PP7_11_net, CLK => Clock, Q => DF1_7_Q);
    DF1_87 : DF1
      port map(D => E_2_net, CLK => Clock, Q => DF1_87_Q);
    BUF_5 : BUFF
      port map(A => DataA(7), Y => BUF_5_Y);
    DF1_144 : DF1
      port map(D => PP3_4_net, CLK => Clock, Q => DF1_144_Q);
    DF1_108 : DF1
      port map(D => E_3_net, CLK => Clock, Q => DF1_108_Q);
    HA1_14 : HA1
      port map(A => DF1_126_Q, B => DF1_38_Q, CO => HA1_14_CO, 
        S => HA1_14_S);
    DF1_14 : DF1
      port map(D => PP7_5_net, CLK => Clock, Q => DF1_14_Q);
    DF1_68 : DF1
      port map(D => PP5_15_net, CLK => Clock, Q => DF1_68_Q);
    OR3_2 : OR3
      port map(A => DataB(1), B => DataB(2), C => DataB(3), Y => 
        OR3_2_Y);
    BUF_30 : BUFF
      port map(A => DataB(5), Y => BUF_30_Y);
    ADD1_Mult_18_inst : ADD1
      port map(A => SumA_17_net, B => SumB_17_net, FCI => 
        ADD1_Mult_17_FCO, S => Mult(18), FCO => ADD1_Mult_18_FCO);
    XOR2_PP2_8_inst : XOR2
      port map(A => AO6_47_Y, B => BUF_34_Y, Y => PP2_8_net);
    XOR2_7 : XOR2
      port map(A => BUF_40_Y, B => DataB(13), Y => XOR2_7_Y);
    DF1_115 : DF1
      port map(D => PP2_12_net, CLK => Clock, Q => DF1_115_Q);
    BUF_0 : BUFF
      port map(A => DataA(14), Y => BUF_0_Y);
    DF1_34 : DF1
      port map(D => PP2_1_net, CLK => Clock, Q => DF1_34_Q);
    FA1_2 : FA1
      port map(A => FA1_17_CO, B => FA1_56_S, CI => FA1_49_S, 
        CO => FA1_2_CO, S => FA1_2_S);
    FA1_20 : FA1
      port map(A => FA1_33_CO, B => FA1_40_CO, CI => FA1_61_S, 
        CO => FA1_20_CO, S => FA1_20_S);
    DF1_132 : DF1
      port map(D => PP5_1_net, CLK => Clock, Q => DF1_132_Q);
    AO6_95 : AO6
      port map(A => BUF_32_Y, B => AO16_6_Y, C => BUF_31_Y, D => 
        XOR2_18_Y, Y => AO6_95_Y);
    BUF_32 : BUFF
      port map(A => DataA(13), Y => BUF_32_Y);
    AO6_40 : AO6
      port map(A => BUF_13_Y, B => AO16_5_Y, C => BUF_44_Y, D => 
        XOR2_8_Y, Y => AO6_40_Y);
    XOR2_23 : XOR2
      port map(A => DataB(3), B => DataB(4), Y => XOR2_23_Y);
    XOR2_PP5_2_inst : XOR2
      port map(A => AO6_72_Y, B => BUF_47_Y, Y => PP5_2_net);
    AO6_26 : AO6
      port map(A => BUF_44_Y, B => AO16_1_Y, C => BUF_19_Y, D => 
        XOR2_10_Y, Y => AO6_26_Y);
    DF1_SumA_23_inst : DF1
      port map(D => FA1_16_CO, CLK => Clock, Q => SumA_23_net);
    XOR2_PP2_15_inst : XOR2
      port map(A => AO6_79_Y, B => BUF_30_Y, Y => PP2_15_net);
    XOR2_29 : XOR2
      port map(A => DataB(9), B => DataB(10), Y => XOR2_29_Y);
    FA1_56 : FA1
      port map(A => FA1_6_CO, B => DF1_39_Q, CI => FA1_55_S, 
        CO => FA1_56_CO, S => FA1_56_S);
    DF1_102 : DF1
      port map(D => PP0_10_net, CLK => Clock, Q => DF1_102_Q);
    DF1_SumA_10_inst : DF1
      port map(D => FA1_23_CO, CLK => Clock, Q => SumA_10_net);
    XOR2_PP3_5_inst : XOR2
      port map(A => AO6_62_Y, B => BUF_12_Y, Y => PP3_5_net);
    XOR2_PP0_9_inst : XOR2
      port map(A => AO6_41_Y, B => BUF_23_Y, Y => PP0_9_net);
    XOR2_PP2_6_inst : XOR2
      port map(A => AO6_9_Y, B => BUF_34_Y, Y => PP2_6_net);
    FA1_54 : FA1
      port map(A => FA1_5_CO, B => FA1_12_CO, CI => FA1_38_S, 
        CO => FA1_54_CO, S => FA1_54_S);
    DF1_152 : DF1
      port map(D => PP7_1_net, CLK => Clock, Q => DF1_152_Q);
    DF1_SumA_15_inst : DF1
      port map(D => FA1_95_CO, CLK => Clock, Q => SumA_15_net);
    XOR2_27 : XOR2
      port map(A => AND2_2_Y, B => BUF_18_Y, Y => XOR2_27_Y);
    DF1_SumA_3_inst : DF1
      port map(D => HA1_3_CO, CLK => Clock, Q => SumA_3_net);
    XOR2_6 : XOR2
      port map(A => DataB(9), B => DataB(10), Y => XOR2_6_Y);
    BUF_7 : BUFF
      port map(A => DataA(6), Y => BUF_7_Y);
    FCINIT_BUFF_0 : FCINIT_BUFF
      port map(A => GND_1_net, FCO => FCINIT_BUFF_0_FCO);
    AO6_36 : AO6
      port map(A => BUF_4_Y, B => AO16_4_Y, C => BUF_2_Y, D => 
        XOR2_29_Y, Y => AO6_36_Y);
    BUF_4 : BUFF
      port map(A => DataA(3), Y => BUF_4_Y);
    FA1_3 : FA1
      port map(A => DF1_48_Q, B => DF1_87_Q, CI => DF1_31_Q, 
        CO => FA1_3_CO, S => FA1_3_S);
    BUF_18 : BUFF
      port map(A => DataB(3), Y => BUF_18_Y);
    FA1_30 : FA1
      port map(A => DF1_78_Q, B => DF1_97_Q, CI => DF1_145_Q, 
        CO => FA1_30_CO, S => FA1_30_S);
    DF1_123 : DF1
      port map(D => PP1_11_net, CLK => Clock, Q => DF1_123_Q);
    BUF_28 : BUFF
      port map(A => DataA(3), Y => BUF_28_Y);
    DF1_89 : DF1
      port map(D => PP7_14_net, CLK => Clock, Q => DF1_89_Q);
    MX2_PP0_16_inst : MX2
      port map(A => MX2_2_Y, B => EBAR, S => AND2A_1_Y, Y => 
        PP0_16_net);
    AO6_9 : AO6
      port map(A => BUF_45_Y, B => AO16_10_Y, C => BUF_7_Y, D => 
        XOR2_21_Y, Y => AO6_9_Y);
    DF1_18 : DF1
      port map(D => PP0_6_net, CLK => Clock, Q => DF1_18_Q);
    DF1_SumB_30_inst : DF1
      port map(D => HA1_4_CO, CLK => Clock, Q => SumB_30_net);
    DF1_SumB_22_inst : DF1
      port map(D => FA1_16_S, CLK => Clock, Q => SumB_22_net);
    AO6_45 : AO6
      port map(A => BUF_21_Y, B => AND2A_0_Y, C => BUF_27_Y, D => 
        DataB(0), Y => AO6_45_Y);
    AO6_13 : AO6
      port map(A => BUF_9_Y, B => AO16_2_Y, C => BUF_15_Y, D => 
        XOR2_6_Y, Y => AO6_13_Y);
    AO6_50 : AO6
      port map(A => BUF_2_Y, B => AO16_4_Y, C => BUF_36_Y, D => 
        XOR2_29_Y, Y => AO6_50_Y);
    DF1_54 : DF1
      port map(D => PP6_6_net, CLK => Clock, Q => DF1_54_Q);
    AND2A_1 : AND2A
      port map(A => DataB(0), B => BUF_23_Y, Y => AND2A_1_Y);
    XOR2_PP6_5_inst : XOR2
      port map(A => AO6_67_Y, B => BUF_17_Y, Y => PP6_5_net);
    XOR2_PP6_8_inst : XOR2
      port map(A => AO6_90_Y, B => BUF_17_Y, Y => PP6_8_net);
    DF1_26 : DF1
      port map(D => PP7_15_net, CLK => Clock, Q => DF1_26_Q);
    DF1_38 : DF1
      port map(D => PP6_12_net, CLK => Clock, Q => DF1_38_Q);
    XOR2_PP4_13_inst : XOR2
      port map(A => AO6_53_Y, B => BUF_33_Y, Y => PP4_13_net);
    XOR2_PP4_3_inst : XOR2
      port map(A => AO6_112_Y, B => BUF_37_Y, Y => PP4_3_net);
    ADD1_Mult_9_inst : ADD1
      port map(A => SumA_8_net, B => SumB_8_net, FCI => 
        ADD1_Mult_8_FCO, S => Mult(9), FCO => ADD1_Mult_9_FCO);
    BUF_10 : BUFF
      port map(A => DataA(9), Y => BUF_10_Y);
    AO6_12 : AO6
      port map(A => BUF_10_Y, B => AO16_7_Y, C => BUF_43_Y, D => 
        XOR2_28_Y, Y => AO6_12_Y);
    FA1_6 : FA1
      port map(A => DF1_67_Q, B => DF1_128_Q, CI => DF1_44_Q, 
        CO => FA1_6_CO, S => FA1_6_S);
    ADD1_Mult_5_inst : ADD1
      port map(A => SumA_4_net, B => SumB_4_net, FCI => 
        ADD1_Mult_4_FCO, S => Mult(5), FCO => ADD1_Mult_5_FCO);
    FA1_60 : FA1
      port map(A => FA1_10_CO, B => HA1_2_CO, CI => FA1_6_S, 
        CO => FA1_60_CO, S => FA1_60_S);
    BUF_20 : BUFF
      port map(A => DataB(15), Y => BUF_20_Y);
    XOR2_PP7_15_inst : XOR2
      port map(A => AO6_69_Y, B => BUF_20_Y, Y => PP7_15_net);
    DF1_SumB_11_inst : DF1
      port map(D => FA1_76_S, CLK => Clock, Q => SumB_11_net);
    XOR2_PP6_9_inst : XOR2
      port map(A => AO6_54_Y, B => BUF_6_Y, Y => PP6_9_net);
    XOR2_PP1_2_inst : XOR2
      port map(A => AO6_29_Y, B => BUF_18_Y, Y => PP1_2_net);
    HA1_15 : HA1
      port map(A => DF1_6_Q, B => DF1_107_Q, CO => HA1_15_CO, 
        S => HA1_15_S);
    BUF_12 : BUFF
      port map(A => DataB(7), Y => BUF_12_Y);
    AOI1_E_0_inst : AOI1
      port map(A => XOR2_26_Y, B => OR3_1_Y, C => AND3_1_Y, Y => 
        E_0_net);
    XOR2_PP1_10_inst : XOR2
      port map(A => AO6_22_Y, B => BUF_11_Y, Y => PP1_10_net);
    XOR2_PP3_15_inst : XOR2
      port map(A => AO6_15_Y, B => BUF_3_Y, Y => PP3_15_net);
    MX2_PP5_16_inst : MX2
      port map(A => MX2_3_Y, B => AO1_4_Y, S => AO16_2_Y, Y => 
        PP5_16_net);
    BUF_22 : BUFF
      port map(A => DataB(15), Y => BUF_22_Y);
    AO6_4 : AO6
      port map(A => BUF_27_Y, B => AND2A_0_Y, C => BUF_28_Y, D => 
        DataB(0), Y => AO6_4_Y);
    BUF_31 : BUFF
      port map(A => DataA(14), Y => BUF_31_Y);
    AO6_55 : AO6
      port map(A => BUF_25_Y, B => AO16_5_Y, C => BUF_4_Y, D => 
        XOR2_8_Y, Y => AO6_55_Y);
    XOR2_PP5_9_inst : XOR2
      port map(A => AO6_82_Y, B => BUF_41_Y, Y => PP5_9_net);
    AO6_114 : AO6
      port map(A => BUF_29_Y, B => AND2A_0_Y, C => BUF_21_Y, D => 
        DataB(0), Y => AO6_114_Y);
    DF1_66 : DF1
      port map(D => PP2_13_net, CLK => Clock, Q => DF1_66_Q);
    XOR2_0 : XOR2
      port map(A => AND2_4_Y, B => BUF_37_Y, Y => XOR2_0_Y);
    DF1_SumA_9_inst : DF1
      port map(D => FA1_64_CO, CLK => Clock, Q => SumA_9_net);
    HA1_S_5_inst : HA1
      port map(A => XOR2_24_Y, B => DataB(11), CO => S_5_net, 
        S => PP5_0_net);
    AO6_94 : AO6
      port map(A => BUF_32_Y, B => AO16_0_Y, C => BUF_31_Y, D => 
        XOR2_5_Y, Y => AO6_94_Y);
    AO6_116 : AO6
      port map(A => BUF_14_Y, B => AO16_9_Y, C => BUF_10_Y, D => 
        XOR2_23_Y, Y => AO6_116_Y);
    DF1_73 : DF1
      port map(D => PP0_15_net, CLK => Clock, Q => DF1_73_Q);
    XOR2_PP6_12_inst : XOR2
      port map(A => AO6_3_Y, B => BUF_6_Y, Y => PP6_12_net);
    DF1_58 : DF1
      port map(D => PP4_0_net, CLK => Clock, Q => DF1_58_Q);
    XOR2_PP0_1_inst : XOR2
      port map(A => AO6_114_Y, B => BUF_26_Y, Y => PP0_1_net);
    XOR2_PP4_1_inst : XOR2
      port map(A => AO6_10_Y, B => BUF_37_Y, Y => PP4_1_net);
    XOR2_PP5_3_inst : XOR2
      port map(A => AO6_52_Y, B => BUF_47_Y, Y => PP5_3_net);
    FA1_55 : FA1
      port map(A => DF1_59_Q, B => DF1_10_Q, CI => DF1_19_Q, 
        CO => FA1_55_CO, S => FA1_55_S);
    DF1_70 : DF1
      port map(D => PP1_12_net, CLK => Clock, Q => DF1_70_Q);
    AO6_105 : AO6
      port map(A => BUF_45_Y, B => AO16_13_Y, C => BUF_7_Y, D => 
        XOR2_25_Y, Y => AO6_105_Y);
    AOI1_E_2_inst : AOI1
      port map(A => XOR2_22_Y, B => OR3_6_Y, C => AND3_2_Y, Y => 
        E_2_net);
    AO6_5 : AO6
      port map(A => BUF_24_Y, B => AO16_9_Y, C => BUF_16_Y, D => 
        XOR2_23_Y, Y => AO6_5_Y);
    DF1_75 : DF1
      port map(D => E_4_net, CLK => Clock, Q => DF1_75_Q);
    DF1_SumB_20_inst : DF1
      port map(D => FA1_53_S, CLK => Clock, Q => SumB_20_net);
    DF1_21 : DF1
      port map(D => S_1_net, CLK => Clock, Q => DF1_21_Q);
    DF1_94 : DF1
      port map(D => PP1_16_net, CLK => Clock, Q => DF1_94_Q);
    AO6_99 : AO6
      port map(A => BUF_43_Y, B => AO16_7_Y, C => BUF_42_Y, D => 
        XOR2_28_Y, Y => AO6_99_Y);
    DF1_SumA_19_inst : DF1
      port map(D => FA1_79_CO, CLK => Clock, Q => SumA_19_net);
    DF1_27 : DF1
      port map(D => PP2_11_net, CLK => Clock, Q => DF1_27_Q);
    DF1_141 : DF1
      port map(D => PP4_4_net, CLK => Clock, Q => DF1_141_Q);
    DF1_SumA_26_inst : DF1
      port map(D => FA1_39_CO, CLK => Clock, Q => SumA_26_net);
    ADD1_Mult_7_inst : ADD1
      port map(A => SumA_6_net, B => SumB_6_net, FCI => 
        ADD1_Mult_6_FCO, S => Mult(7), FCO => ADD1_Mult_7_FCO);
    DF1_42 : DF1
      port map(D => PP1_3_net, CLK => Clock, Q => DF1_42_Q);
    AO6_44 : AO6
      port map(A => BUF_36_Y, B => AO16_5_Y, C => BUF_13_Y, D => 
        XOR2_8_Y, Y => AO6_44_Y);
    DF1_SumB_25_inst : DF1
      port map(D => FA1_39_S, CLK => Clock, Q => SumB_25_net);
    AOI1_E_7_inst : AOI1
      port map(A => XOR2_11_Y, B => OR3_4_Y, C => AND3_7_Y, Y => 
        E_7_net);
    XOR2_21 : XOR2
      port map(A => DataB(3), B => DataB(4), Y => XOR2_21_Y);
    AO6_17 : AO6
      port map(A => BUF_42_Y, B => AO16_9_Y, C => BUF_24_Y, D => 
        XOR2_23_Y, Y => AO6_17_Y);
    XOR2_PP0_2_inst : XOR2
      port map(A => AO6_45_Y, B => BUF_26_Y, Y => PP0_2_net);
    XOR2_PP6_3_inst : XOR2
      port map(A => AO6_55_Y, B => BUF_17_Y, Y => PP6_3_net);
    DF1_16 : DF1
      port map(D => PP6_0_net, CLK => Clock, Q => DF1_16_Q);
    DF1_148 : DF1
      port map(D => S_2_net, CLK => Clock, Q => DF1_148_Q);
    DF1_SumA_28_inst : DF1
      port map(D => FA1_19_CO, CLK => Clock, Q => SumA_28_net);
    XOR2_PP0_11_inst : XOR2
      port map(A => AO6_92_Y, B => BUF_23_Y, Y => PP0_11_net);
    XOR2_14 : XOR2
      port map(A => AND2_5_Y, B => BUF_12_Y, Y => XOR2_14_Y);
    AO1_EBAR : AO1
      port map(A => XOR2_26_Y, B => OR3_1_Y, C => AND3_1_Y, Y => 
        EBAR);
    BUF_11 : BUFF
      port map(A => DataB(3), Y => BUF_11_Y);
    DF1_119 : DF1
      port map(D => PP5_12_net, CLK => Clock, Q => DF1_119_Q);
    BUF_21 : BUFF
      port map(A => DataA(1), Y => BUF_21_Y);
    FA1_79 : FA1
      port map(A => FA1_20_CO, B => FA1_60_S, CI => FA1_17_S, 
        CO => FA1_79_CO, S => FA1_79_S);
    DF1_36 : DF1
      port map(D => PP1_1_net, CLK => Clock, Q => DF1_36_Q);
    FA1_92 : FA1
      port map(A => FA1_1_CO, B => FA1_68_CO, CI => FA1_22_S, 
        CO => FA1_92_CO, S => FA1_92_S);
    AO6_18 : AO6
      port map(A => BUF_27_Y, B => AO16_11_Y, C => BUF_28_Y, D => 
        XOR2_17_Y, Y => AO6_18_Y);
    DF1_61 : DF1
      port map(D => PP1_10_net, CLK => Clock, Q => DF1_61_Q);
    XOR2_PP5_11_inst : XOR2
      port map(A => AO6_13_Y, B => BUF_41_Y, Y => PP5_11_net);
    XOR2_4 : XOR2
      port map(A => DataB(1), B => DataB(2), Y => XOR2_4_Y);
    AO6_49 : AO6
      port map(A => BUF_19_Y, B => AO16_0_Y, C => BUF_38_Y, D => 
        XOR2_5_Y, Y => AO6_49_Y);
    DF1_SumA_13_inst : DF1
      port map(D => FA1_73_CO, CLK => Clock, Q => SumA_13_net);
    XOR2_PP1_9_inst : XOR2
      port map(A => AO6_1_Y, B => BUF_11_Y, Y => PP1_9_net);
    DF1_67 : DF1
      port map(D => PP3_13_net, CLK => Clock, Q => DF1_67_Q);
    AO6_0 : AO6
      port map(A => BUF_4_Y, B => AO16_5_Y, C => BUF_2_Y, D => 
        XOR2_8_Y, Y => AO6_0_Y);
    BUF_47 : BUFF
      port map(A => DataB(11), Y => BUF_47_Y);
    HA1_1 : HA1
      port map(A => DF1_14_Q, B => DF1_53_Q, CO => HA1_1_CO, S => 
        HA1_1_S);
    HA1_10 : HA1
      port map(A => DF1_118_Q, B => VCC_1_net, CO => HA1_10_CO, 
        S => HA1_10_S);
    XOR2_PP5_6_inst : XOR2
      port map(A => AO6_25_Y, B => BUF_47_Y, Y => PP5_6_net);
    AO6_54 : AO6
      port map(A => BUF_19_Y, B => AO16_8_Y, C => BUF_38_Y, D => 
        XOR2_3_Y, Y => AO6_54_Y);
    DF1_136 : DF1
      port map(D => PP5_8_net, CLK => Clock, Q => DF1_136_Q);
    XOR2_PP0_14_inst : XOR2
      port map(A => AO6_30_Y, B => BUF_23_Y, Y => PP0_14_net);
    ADD1_Mult_4_inst : ADD1
      port map(A => SumA_3_net, B => SumB_3_net, FCI => 
        ADD1_Mult_3_FCO, S => Mult(4), FCO => ADD1_Mult_4_FCO);
    DF1_142 : DF1
      port map(D => S_3_net, CLK => Clock, Q => DF1_142_Q);
    DF1_98 : DF1
      port map(D => PP3_7_net, CLK => Clock, Q => DF1_98_Q);
    DF1_SumA_8_inst : DF1
      port map(D => FA1_80_CO, CLK => Clock, Q => SumA_8_net);
    AO6_110 : AO6
      port map(A => BUF_7_Y, B => AO16_11_Y, C => BUF_5_Y, D => 
        XOR2_17_Y, Y => AO6_110_Y);
    AND2_1 : AND2
      port map(A => XOR2_21_Y, B => BUF_29_Y, Y => AND2_1_Y);
    OR3_3 : OR3
      port map(A => DataB(9), B => DataB(10), C => DataB(11), 
        Y => OR3_3_Y);
    DF1_29 : DF1
      port map(D => S_7_net, CLK => Clock, Q => DF1_29_Q);
    DF1_SumB_14_inst : DF1
      port map(D => FA1_95_S, CLK => Clock, Q => SumB_14_net);
    DF1_SumB_2_inst : DF1
      port map(D => HA1_3_S, CLK => Clock, Q => SumB_2_net);
    XOR2_PP4_12_inst : XOR2
      port map(A => AO6_37_Y, B => BUF_33_Y, Y => PP4_12_net);
    HA1_S_4_inst : HA1
      port map(A => XOR2_0_Y, B => DataB(9), CO => S_4_net, S => 
        PP4_0_net);
    DF1_106 : DF1
      port map(D => PP3_14_net, CLK => Clock, Q => DF1_106_Q);
    AND2_7 : AND2
      port map(A => XOR2_2_Y, B => BUF_8_Y, Y => AND2_7_Y);
    XOR2_PP5_14_inst : XOR2
      port map(A => AO6_115_Y, B => BUF_41_Y, Y => PP5_14_net);
    BUF_33 : BUFF
      port map(A => DataB(9), Y => BUF_33_Y);
    AO6_73 : AO6
      port map(A => BUF_28_Y, B => AND2A_0_Y, C => BUF_39_Y, D => 
        DataB(0), Y => AO6_73_Y);
    XOR2_PP0_6_inst : XOR2
      port map(A => AO6_76_Y, B => BUF_26_Y, Y => PP0_6_net);
    XOR2_PP3_1_inst : XOR2
      port map(A => AO6_16_Y, B => BUF_12_Y, Y => PP3_1_net);
    XOR2_15 : XOR2
      port map(A => BUF_46_Y, B => DataB(7), Y => XOR2_15_Y);
    HA1_6 : HA1
      port map(A => DF1_52_Q, B => DF1_60_Q, CO => HA1_6_CO, S => 
        HA1_6_S);
    FCEND_BUFF_0 : FCEND_BUFF
      port map(FCI => ADD1_Mult_31_FCO, CO => FCEND_BUFF_0_CO);
    AO6_111 : AO6
      port map(A => BUF_2_Y, B => AO16_12_Y, C => BUF_36_Y, D => 
        XOR2_2_Y, Y => AO6_111_Y);
    FA1_19 : FA1
      port map(A => HA1_5_S, B => DF1_89_Q, CI => FA1_65_CO, 
        CO => FA1_19_CO, S => FA1_19_S);
    MX2_4 : MX2
      port map(A => BUF_20_Y, B => XOR2_11_Y, S => XOR2_18_Y, 
        Y => MX2_4_Y);
    AO6_59 : AO6
      port map(A => BUF_24_Y, B => AO16_7_Y, C => BUF_16_Y, D => 
        XOR2_28_Y, Y => AO6_59_Y);
    AO6_60 : AO6
      port map(A => BUF_44_Y, B => AO16_4_Y, C => BUF_19_Y, D => 
        XOR2_29_Y, Y => AO6_60_Y);
    DF1_56 : DF1
      port map(D => PP6_13_net, CLK => Clock, Q => DF1_56_Q);
    FA1_5 : FA1
      port map(A => DF1_82_Q, B => DF1_33_Q, CI => HA1_13_CO, 
        CO => FA1_5_CO, S => FA1_5_S);
    AND3_4 : AND3
      port map(A => DataB(5), B => DataB(6), C => DataB(7), Y => 
        AND3_4_Y);
    XOR2_PP2_2_inst : XOR2
      port map(A => AO6_106_Y, B => BUF_34_Y, Y => PP2_2_net);
    AO6_72 : AO6
      port map(A => BUF_35_Y, B => AO16_4_Y, C => BUF_25_Y, D => 
        XOR2_29_Y, Y => AO6_72_Y);
    FA1_50 : FA1
      port map(A => DF1_5_Q, B => VCC_1_net, CI => DF1_129_Q, 
        CO => FA1_50_CO, S => FA1_50_S);
    AO6_83 : AO6
      port map(A => BUF_4_Y, B => AO16_1_Y, C => BUF_2_Y, D => 
        XOR2_10_Y, Y => AO6_83_Y);
    DF1_114 : DF1
      port map(D => PP0_1_net, CLK => Clock, Q => DF1_114_Q);
    DF1_11 : DF1
      port map(D => PP3_12_net, CLK => Clock, Q => DF1_11_Q);
    BUF_8 : BUFF
      port map(A => DataA(0), Y => BUF_8_Y);
    AO6_96 : AO6
      port map(A => BUF_25_Y, B => AO16_12_Y, C => BUF_4_Y, D => 
        XOR2_2_Y, Y => AO6_96_Y);
    HA1_3 : HA1
      port map(A => DF1_36_Q, B => DF1_111_Q, CO => HA1_3_CO, 
        S => HA1_3_S);
    DF1_17 : DF1
      port map(D => PP2_7_net, CLK => Clock, Q => DF1_17_Q);
    AOI1_E_4_inst : AOI1
      port map(A => XOR2_20_Y, B => OR3_7_Y, C => AND3_0_Y, Y => 
        E_4_net);
    DF1_69 : DF1
      port map(D => PP6_9_net, CLK => Clock, Q => DF1_69_Q);
    AO6_82 : AO6
      port map(A => BUF_19_Y, B => AO16_2_Y, C => BUF_38_Y, D => 
        XOR2_6_Y, Y => AO6_82_Y);
    AND3_1 : AND3
      port map(A => GND_1_net, B => DataB(0), C => DataB(1), Y => 
        AND3_1_Y);
    XOR2_22 : XOR2
      port map(A => BUF_46_Y, B => DataB(5), Y => XOR2_22_Y);
    DF1_31 : DF1
      port map(D => PP4_13_net, CLK => Clock, Q => DF1_31_Q);
    FA1_49 : FA1
      port map(A => FA1_60_CO, B => FA1_11_CO, CI => FA1_27_S, 
        CO => FA1_49_CO, S => FA1_49_S);
    DF1_SumB_29_inst : DF1
      port map(D => FA1_88_CO, CLK => Clock, Q => SumB_29_net);
    AO16_13 : AO16
      port map(A => DataB(1), B => DataB(2), C => BUF_18_Y, Y => 
        AO16_13_Y);
    DF1_127 : DF1
      port map(D => PP3_0_net, CLK => Clock, Q => DF1_127_Q);
    DF1_37 : DF1
      port map(D => PP4_10_net, CLK => Clock, Q => DF1_37_Q);
    XOR2_PP6_1_inst : XOR2
      port map(A => AO6_97_Y, B => BUF_17_Y, Y => PP6_1_net);
    AO6_119 : AO6
      port map(A => BUF_10_Y, B => AO16_9_Y, C => BUF_43_Y, D => 
        XOR2_23_Y, Y => AO6_119_Y);
    FA1_89 : FA1
      port map(A => DF1_64_Q, B => DF1_17_Q, CI => DF1_149_Q, 
        CO => FA1_89_CO, S => FA1_89_S);
    XOR2_10 : XOR2
      port map(A => DataB(7), B => DataB(8), Y => XOR2_10_Y);
    XOR2_PP3_6_inst : XOR2
      port map(A => AO6_103_Y, B => BUF_12_Y, Y => PP3_6_net);
    AO6_65 : AO6
      port map(A => BUF_8_Y, B => AO16_4_Y, C => BUF_35_Y, D => 
        XOR2_29_Y, Y => AO6_65_Y);
    XOR2_PP1_13_inst : XOR2
      port map(A => AO6_113_Y, B => BUF_11_Y, Y => PP1_13_net);
    ADD1_Mult_22_inst : ADD1
      port map(A => SumA_21_net, B => SumB_21_net, FCI => 
        ADD1_Mult_21_FCO, S => Mult(22), FCO => ADD1_Mult_22_FCO);
    XOR2_26 : XOR2
      port map(A => BUF_46_Y, B => DataB(1), Y => XOR2_26_Y);
    HA1_S_7_inst : HA1
      port map(A => XOR2_12_Y, B => DataB(15), CO => S_7_net, 
        S => PP7_0_net);
    AO6_23 : AO6
      port map(A => BUF_0_Y, B => AO16_3_Y, C => BUF_46_Y, D => 
        XOR2_4_Y, Y => AO6_23_Y);
    XOR2_PP2_1_inst : XOR2
      port map(A => AO6_24_Y, B => BUF_34_Y, Y => PP2_1_net);
    AO6_46 : AO6
      port map(A => BUF_28_Y, B => AO16_13_Y, C => BUF_39_Y, D => 
        XOR2_25_Y, Y => AO6_46_Y);
    XOR2_PP2_10_inst : XOR2
      port map(A => AO6_119_Y, B => BUF_30_Y, Y => PP2_10_net);
    BUF_13 : BUFF
      port map(A => DataA(6), Y => BUF_13_Y);
    DF1_120 : DF1
      port map(D => PP1_0_net, CLK => Clock, Q => DF1_120_Q);
    FA1_29 : FA1
      port map(A => DF1_135_Q, B => DF1_90_Q, CI => DF1_88_Q, 
        CO => FA1_29_CO, S => FA1_29_S);
    AO6_11 : AO6
      port map(A => BUF_42_Y, B => AND2A_1_Y, C => BUF_24_Y, D => 
        DataB(0), Y => AO6_11_Y);
    AND2_3 : AND2
      port map(A => XOR2_8_Y, B => BUF_8_Y, Y => AND2_3_Y);
    BUF_23 : BUFF
      port map(A => DataB(1), Y => BUF_23_Y);
    XOR2_PP1_6_inst : XOR2
      port map(A => AO6_105_Y, B => BUF_18_Y, Y => PP1_6_net);
    FA1_78 : FA1
      port map(A => FA1_45_CO, B => FA1_50_S, CI => FA1_70_S, 
        CO => FA1_78_CO, S => FA1_78_S);
    DF1_SumB_23_inst : DF1
      port map(D => FA1_78_S, CLK => Clock, Q => SumB_23_net);
    FA1_72 : FA1
      port map(A => FA1_58_CO, B => FA1_89_S, CI => FA1_57_S, 
        CO => FA1_72_CO, S => FA1_72_S);
    XOR2_PP7_3_inst : XOR2
      port map(A => AO6_96_Y, B => BUF_22_Y, Y => PP7_3_net);
    AO6_22 : AO6
      port map(A => BUF_10_Y, B => AO16_3_Y, C => BUF_43_Y, D => 
        XOR2_4_Y, Y => AO6_22_Y);
    MX2_PP7_16_inst : MX2
      port map(A => MX2_4_Y, B => AO1_3_Y, S => AO16_6_Y, Y => 
        PP7_16_net);
    DF1_74 : DF1
      port map(D => PP4_7_net, CLK => Clock, Q => DF1_74_Q);
    DF1_82 : DF1
      port map(D => PP5_2_net, CLK => Clock, Q => DF1_82_Q);
    DF1_51 : DF1
      port map(D => PP3_1_net, CLK => Clock, Q => DF1_51_Q);
    BUF_39 : BUFF
      port map(A => DataA(4), Y => BUF_39_Y);
    XOR2_PP3_4_inst : XOR2
      port map(A => AO6_43_Y, B => BUF_12_Y, Y => PP3_4_net);
    AO6_6 : AO6
      port map(A => BUF_19_Y, B => AO16_6_Y, C => BUF_38_Y, D => 
        XOR2_18_Y, Y => AO6_6_Y);
    DF1_4 : DF1
      port map(D => PP6_16_net, CLK => Clock, Q => DF1_4_Q);
    DF1_19 : DF1
      port map(D => PP6_8_net, CLK => Clock, Q => DF1_19_Q);
    AO6_33 : AO6
      port map(A => BUF_42_Y, B => AO16_3_Y, C => BUF_24_Y, D => 
        XOR2_4_Y, Y => AO6_33_Y);
    DF1_96 : DF1
      port map(D => PP3_10_net, CLK => Clock, Q => DF1_96_Q);
    DF1_57 : DF1
      port map(D => PP7_12_net, CLK => Clock, Q => DF1_57_Q);
    DF1_SumA_16_inst : DF1
      port map(D => FA1_59_CO, CLK => Clock, Q => SumA_16_net);
    AO6_77 : AO6
      port map(A => BUF_28_Y, B => AO16_10_Y, C => BUF_39_Y, D => 
        XOR2_21_Y, Y => AO6_77_Y);
    AND2A_0 : AND2A
      port map(A => DataB(0), B => BUF_26_Y, Y => AND2A_0_Y);
    DF1_39 : DF1
      port map(D => PP7_6_net, CLK => Clock, Q => DF1_39_Q);
    DF1_SumA_1_inst : DF1
      port map(D => DF1_25_Q, CLK => Clock, Q => SumA_1_net);
    DF1_125 : DF1
      port map(D => PP2_2_net, CLK => Clock, Q => DF1_125_Q);
    XOR2_PP4_8_inst : XOR2
      port map(A => AO6_26_Y, B => BUF_37_Y, Y => PP4_8_net);
    AO6_56 : AO6
      port map(A => BUF_38_Y, B => AO16_8_Y, C => BUF_9_Y, D => 
        XOR2_3_Y, Y => AO6_56_Y);
    FA1_39 : FA1
      port map(A => FA1_52_CO, B => FA1_47_CO, CI => FA1_8_S, 
        CO => FA1_39_CO, S => FA1_39_S);
    AO6_32 : AO6
      port map(A => BUF_39_Y, B => AND2A_0_Y, C => BUF_45_Y, D => 
        DataB(0), Y => AO6_32_Y);
    DF1_SumA_21_inst : DF1
      port map(D => FA1_53_CO, CLK => Clock, Q => SumA_21_net);
    ADD1_Mult_25_inst : ADD1
      port map(A => SumA_24_net, B => SumB_24_net, FCI => 
        ADD1_Mult_24_FCO, S => Mult(25), FCO => ADD1_Mult_25_FCO);
    AO16_8 : AO16
      port map(A => DataB(11), B => DataB(12), C => BUF_6_Y, Y => 
        AO16_8_Y);
    DF1_SumA_18_inst : DF1
      port map(D => FA1_4_CO, CLK => Clock, Q => SumA_18_net);
    AO6_78 : AO6
      port map(A => BUF_16_Y, B => AO16_3_Y, C => BUF_0_Y, D => 
        XOR2_4_Y, Y => AO6_78_Y);
    DF1_133 : DF1
      port map(D => PP2_14_net, CLK => Clock, Q => DF1_133_Q);
    AO6_87 : AO6
      port map(A => BUF_9_Y, B => AO16_0_Y, C => BUF_15_Y, D => 
        XOR2_5_Y, Y => AO6_87_Y);
    XOR2_13 : XOR2
      port map(A => BUF_46_Y, B => DataB(3), Y => XOR2_13_Y);
    XOR2_2 : XOR2
      port map(A => DataB(13), B => DataB(14), Y => XOR2_2_Y);
    XOR2_3 : XOR2
      port map(A => DataB(11), B => DataB(12), Y => XOR2_3_Y);
    FA1_18 : FA1
      port map(A => DF1_113_Q, B => DF1_100_Q, CI => HA1_8_S, 
        CO => FA1_18_CO, S => FA1_18_S);
    XOR2_PP7_10_inst : XOR2
      port map(A => AO6_34_Y, B => BUF_20_Y, Y => PP7_10_net);
    FA1_12 : FA1
      port map(A => DF1_16_Q, B => DF1_141_Q, CI => FA1_94_S, 
        CO => FA1_12_CO, S => FA1_12_S);
    XOR2_19 : XOR2
      port map(A => BUF_40_Y, B => DataB(11), Y => XOR2_19_Y);
    HA1_7 : HA1
      port map(A => DF1_79_Q, B => DF1_30_Q, CO => HA1_7_CO, S => 
        HA1_7_S);
    AO1_2 : AO1
      port map(A => XOR2_22_Y, B => OR3_6_Y, C => AND3_2_Y, Y => 
        AO1_2_Y);
    XOR2_PP3_7_inst : XOR2
      port map(A => AO6_110_Y, B => BUF_12_Y, Y => PP3_7_net);
    HA1_S_1_inst : HA1
      port map(A => XOR2_27_Y, B => DataB(3), CO => S_1_net, S => 
        PP1_0_net);
    DF1_103 : DF1
      port map(D => PP4_2_net, CLK => Clock, Q => DF1_103_Q);
    XOR2_PP0_4_inst : XOR2
      port map(A => AO6_73_Y, B => BUF_26_Y, Y => PP0_4_net);
    AO6_88 : AO6
      port map(A => BUF_0_Y, B => AND2A_1_Y, C => BUF_46_Y, D => 
        DataB(0), Y => AO6_88_Y);
    XOR2_PP3_10_inst : XOR2
      port map(A => AO6_12_Y, B => BUF_3_Y, Y => PP3_10_net);
    FA1_69 : FA1
      port map(A => FA1_70_CO, B => FA1_47_S, CI => FA1_52_S, 
        CO => FA1_69_CO, S => FA1_69_S);
    XOR2_PP1_8_inst : XOR2
      port map(A => AO6_98_Y, B => BUF_18_Y, Y => PP1_8_net);
    XOR2_PP7_4_inst : XOR2
      port map(A => AO6_7_Y, B => BUF_22_Y, Y => PP7_4_net);
    BUF_34 : BUFF
      port map(A => DataB(5), Y => BUF_34_Y);
    HA1_2 : HA1
      port map(A => DF1_80_Q, B => DF1_54_Q, CO => HA1_2_CO, S => 
        HA1_2_S);
    DF1_78 : DF1
      port map(D => PP1_6_net, CLK => Clock, Q => DF1_78_Q);
    XOR2_PP3_9_inst : XOR2
      port map(A => AO6_86_Y, B => BUF_3_Y, Y => PP3_9_net);
    XOR2_PP6_11_inst : XOR2
      port map(A => AO6_102_Y, B => BUF_6_Y, Y => PP6_11_net);
    DF1_SumB_9_inst : DF1
      port map(D => FA1_23_S, CLK => Clock, Q => SumB_9_net);
    AO6_64 : AO6
      port map(A => BUF_35_Y, B => AO16_5_Y, C => BUF_25_Y, D => 
        XOR2_8_Y, Y => AO6_64_Y);
    XOR2_17 : XOR2
      port map(A => DataB(5), B => DataB(6), Y => XOR2_17_Y);
    AO6_104 : AO6
      port map(A => BUF_38_Y, B => AO16_2_Y, C => BUF_9_Y, D => 
        XOR2_6_Y, Y => AO6_104_Y);
    XOR2_PP0_15_inst : XOR2
      port map(A => AO6_88_Y, B => BUF_23_Y, Y => PP0_15_net);
    ADD1_Mult_27_inst : ADD1
      port map(A => SumA_26_net, B => SumB_26_net, FCI => 
        ADD1_Mult_26_FCO, S => Mult(27), FCO => ADD1_Mult_27_FCO);
    DF1_59 : DF1
      port map(D => PP4_12_net, CLK => Clock, Q => DF1_59_Q);
    FA1_48 : FA1
      port map(A => FA1_56_CO, B => FA1_27_CO, CI => FA1_68_S, 
        CO => FA1_48_CO, S => FA1_48_S);
    OR3_1 : OR3
      port map(A => GND_1_net, B => DataB(0), C => DataB(1), Y => 
        OR3_1_Y);
    FA1_42 : FA1
      port map(A => DF1_27_Q, B => DF1_73_Q, CI => DF1_74_Q, 
        CO => FA1_42_CO, S => FA1_42_S);
    DF1_SumB_1_inst : DF1
      port map(D => DF1_120_Q, CLK => Clock, Q => SumB_1_net);
    XOR2_PP5_8_inst : XOR2
      port map(A => AO6_60_Y, B => BUF_47_Y, Y => PP5_8_net);
    BUF_19 : BUFF
      port map(A => DataA(8), Y => BUF_19_Y);
    XOR2_PP6_7_inst : XOR2
      port map(A => AO6_40_Y, B => BUF_17_Y, Y => PP6_7_net);
    AO6_106 : AO6
      port map(A => BUF_21_Y, B => AO16_10_Y, C => BUF_27_Y, D => 
        XOR2_21_Y, Y => AO6_106_Y);
    FA1_88 : FA1
      port map(A => DF1_26_Q, B => DF1_65_Q, CI => HA1_5_CO, 
        CO => FA1_88_CO, S => FA1_88_S);
    BUF_45 : BUFF
      port map(A => DataA(5), Y => BUF_45_Y);
    DF1_146 : DF1
      port map(D => PP7_7_net, CLK => Clock, Q => DF1_146_Q);
    FA1_82 : FA1
      port map(A => DF1_148_Q, B => DF1_34_Q, CI => HA1_11_S, 
        CO => FA1_82_CO, S => FA1_82_S);
    DF1_SumB_17_inst : DF1
      port map(D => FA1_4_S, CLK => Clock, Q => SumB_17_net);
    XOR2_PP5_15_inst : XOR2
      port map(A => AO6_57_Y, B => BUF_41_Y, Y => PP5_15_net);
    BUF_29 : BUFF
      port map(A => DataA(0), Y => BUF_29_Y);
    DF1_91 : DF1
      port map(D => PP5_4_net, CLK => Clock, Q => DF1_91_Q);
    AO6_27 : AO6
      port map(A => BUF_39_Y, B => AO16_10_Y, C => BUF_45_Y, D => 
        XOR2_21_Y, Y => AO6_27_Y);
    XOR2_PP1_5_inst : XOR2
      port map(A => AO6_35_Y, B => BUF_18_Y, Y => PP1_5_net);
    XOR2_PP6_14_inst : XOR2
      port map(A => AO6_74_Y, B => BUF_6_Y, Y => PP6_14_net);
    DF1_97 : DF1
      port map(D => PP0_8_net, CLK => Clock, Q => DF1_97_Q);
    DF1_111 : DF1
      port map(D => PP0_3_net, CLK => Clock, Q => DF1_111_Q);
    XOR2_PP1_3_inst : XOR2
      port map(A => AO6_66_Y, B => BUF_18_Y, Y => PP1_3_net);
    XOR2_PP2_5_inst : XOR2
      port map(A => AO6_27_Y, B => BUF_34_Y, Y => PP2_5_net);
    AO6_69 : AO6
      port map(A => BUF_31_Y, B => AO16_6_Y, C => BUF_40_Y, D => 
        XOR2_18_Y, Y => AO6_69_Y);
    XOR2_PP2_7_inst : XOR2
      port map(A => AO6_80_Y, B => BUF_34_Y, Y => PP2_7_net);
    XOR2_PP4_4_inst : XOR2
      port map(A => AO6_83_Y, B => BUF_37_Y, Y => PP4_4_net);
    AO6_28 : AO6
      port map(A => BUF_13_Y, B => AO16_4_Y, C => BUF_44_Y, D => 
        XOR2_29_Y, Y => AO6_28_Y);
    BUF_46 : BUFF
      port map(A => DataA(15), Y => BUF_46_Y);
    FA1_91 : FA1
      port map(A => FA1_8_CO, B => HA1_10_CO, CI => FA1_65_S, 
        CO => FA1_91_CO, S => FA1_91_S);
    AO16_3 : AO16
      port map(A => DataB(1), B => DataB(2), C => BUF_11_Y, Y => 
        AO16_3_Y);
    HA1_S_2_inst : HA1
      port map(A => XOR2_9_Y, B => DataB(5), CO => S_2_net, S => 
        PP2_0_net);
    XOR2_PP2_9_inst : XOR2
      port map(A => AO6_116_Y, B => BUF_30_Y, Y => PP2_9_net);
    FA1_28 : FA1
      port map(A => DF1_49_Q, B => DF1_102_Q, CI => DF1_103_Q, 
        CO => FA1_28_CO, S => FA1_28_S);
    DF1_118 : DF1
      port map(D => PP5_16_net, CLK => Clock, Q => DF1_118_Q);
    FA1_22 : FA1
      port map(A => DF1_9_Q, B => DF1_119_Q, CI => FA1_3_CO, 
        CO => FA1_22_CO, S => FA1_22_S);
    XOR2_PP1_12_inst : XOR2
      port map(A => AO6_33_Y, B => BUF_11_Y, Y => PP1_12_net);
    HA1_S_3_inst : HA1
      port map(A => XOR2_14_Y, B => DataB(7), CO => S_3_net, S => 
        PP3_0_net);
    AO6_37 : AO6
      port map(A => BUF_15_Y, B => AO16_0_Y, C => BUF_1_Y, D => 
        XOR2_5_Y, Y => AO6_37_Y);
    DF1_SumB_26_inst : DF1
      port map(D => FA1_91_S, CLK => Clock, Q => SumB_26_net);
    DF1_Mult_0_inst : DF1
      port map(D => DF1_117_Q, CLK => Clock, Q => Mult(0));
    DF1_SumA_0_inst : DF1
      port map(D => DF1_114_Q, CLK => Clock, Q => SumA_0_net);
    AOI1_E_6_inst : AOI1
      port map(A => XOR2_7_Y, B => OR3_0_Y, C => AND3_3_Y, Y => 
        E_6_net);
    AO6_38 : AO6
      port map(A => BUF_5_Y, B => AND2A_0_Y, C => BUF_14_Y, D => 
        DataB(0), Y => AO6_38_Y);
    BUF_14 : BUFF
      port map(A => DataA(8), Y => BUF_14_Y);
    DF1_SumA_2_inst : DF1
      port map(D => DF1_21_Q, CLK => Clock, Q => SumA_2_net);
    DF1_43 : DF1
      port map(D => PP3_8_net, CLK => Clock, Q => DF1_43_Q);
    AO16_5 : AO16
      port map(A => DataB(11), B => DataB(12), C => BUF_17_Y, 
        Y => AO16_5_Y);
    BUF_24 : BUFF
      port map(A => DataA(12), Y => BUF_24_Y);
    DF1_SumB_28_inst : DF1
      port map(D => FA1_88_S, CLK => Clock, Q => SumB_28_net);
    DF1_112 : DF1
      port map(D => PP1_9_net, CLK => Clock, Q => DF1_112_Q);
    FA1_38 : FA1
      port map(A => HA1_0_S, B => DF1_3_Q, CI => FA1_63_S, CO => 
        FA1_38_CO, S => FA1_38_S);
    DF1_40 : DF1
      port map(D => S_6_net, CLK => Clock, Q => DF1_40_Q);
    FA1_32 : FA1
      port map(A => HA1_15_S, B => DF1_92_Q, CI => FA1_30_CO, 
        CO => FA1_32_CO, S => FA1_32_S);
    AO6_71 : AO6
      port map(A => BUF_2_Y, B => AO16_1_Y, C => BUF_36_Y, D => 
        XOR2_10_Y, Y => AO6_71_Y);
    AO16_0 : AO16
      port map(A => DataB(7), B => DataB(8), C => BUF_33_Y, Y => 
        AO16_0_Y);
    AO1_1 : AO1
      port map(A => XOR2_15_Y, B => OR3_5_Y, C => AND3_4_Y, Y => 
        AO1_1_Y);
    BUF_6 : BUFF
      port map(A => DataB(13), Y => BUF_6_Y);
    XOR2_PP4_11_inst : XOR2
      port map(A => AO6_87_Y, B => BUF_33_Y, Y => PP4_11_net);
    DF1_SumA_24_inst : DF1
      port map(D => FA1_78_CO, CLK => Clock, Q => SumA_24_net);
    XOR2_PP7_1_inst : XOR2
      port map(A => AO6_14_Y, B => BUF_22_Y, Y => PP7_1_net);
    DF1_99 : DF1
      port map(D => PP4_15_net, CLK => Clock, Q => DF1_99_Q);
    BUF_3 : BUFF
      port map(A => DataB(7), Y => BUF_3_Y);
    DF1_22 : DF1
      port map(D => PP5_11_net, CLK => Clock, Q => DF1_22_Q);
    DF1_45 : DF1
      port map(D => PP0_14_net, CLK => Clock, Q => DF1_45_Q);
    DF1_8 : DF1
      port map(D => PP1_4_net, CLK => Clock, Q => DF1_8_Q);
    ADD1_Mult_12_inst : ADD1
      port map(A => SumA_11_net, B => SumB_11_net, FCI => 
        ADD1_Mult_11_FCO, S => Mult(12), FCO => ADD1_Mult_12_FCO);
    MX2_2 : MX2
      port map(A => BUF_23_Y, B => XOR2_26_Y, S => DataB(0), Y => 
        MX2_2_Y);
    XOR2_PP4_9_inst : XOR2
      port map(A => AO6_49_Y, B => BUF_33_Y, Y => PP4_9_net);
    XOR2_PP2_13_inst : XOR2
      port map(A => AO6_5_Y, B => BUF_30_Y, Y => PP2_13_net);
    AO6_81 : AO6
      port map(A => BUF_43_Y, B => AO16_9_Y, C => BUF_42_Y, D => 
        XOR2_23_Y, Y => AO6_81_Y);
    DF1_76 : DF1
      port map(D => PP2_15_net, CLK => Clock, Q => DF1_76_Q);
    AO6_100 : AO6
      port map(A => BUF_42_Y, B => AO16_7_Y, C => BUF_24_Y, D => 
        XOR2_28_Y, Y => AO6_100_Y);
    FA1_68 : FA1
      port map(A => FA1_55_CO, B => DF1_69_Q, CI => FA1_3_S, 
        CO => FA1_68_CO, S => FA1_68_S);
    FA1_62 : FA1
      port map(A => DF1_132_Q, B => DF1_81_Q, CI => HA1_13_S, 
        CO => FA1_62_CO, S => FA1_62_S);
    AO16_9 : AO16
      port map(A => DataB(3), B => DataB(4), C => BUF_30_Y, Y => 
        AO16_9_Y);
    XOR2_11 : XOR2
      port map(A => BUF_40_Y, B => DataB(15), Y => XOR2_11_Y);
    XOR2_PP4_14_inst : XOR2
      port map(A => AO6_94_Y, B => BUF_33_Y, Y => PP4_14_net);
    AO16_12 : AO16
      port map(A => DataB(13), B => DataB(14), C => BUF_22_Y, 
        Y => AO16_12_Y);
    AO6_101 : AO6
      port map(A => BUF_9_Y, B => AO16_6_Y, C => BUF_15_Y, D => 
        XOR2_18_Y, Y => AO6_101_Y);
    XOR2_PP3_3_inst : XOR2
      port map(A => AO6_18_Y, B => BUF_12_Y, Y => PP3_3_net);
    ADD1_Mult_24_inst : ADD1
      port map(A => SumA_23_net, B => SumB_23_net, FCI => 
        ADD1_Mult_23_FCO, S => Mult(24), FCO => ADD1_Mult_24_FCO);
    DF1_129 : DF1
      port map(D => PP5_14_net, CLK => Clock, Q => DF1_129_Q);
    HA1_0 : HA1
      port map(A => DF1_138_Q, B => DF1_98_Q, CO => HA1_0_CO, 
        S => HA1_0_S);
    XOR2_PP3_8_inst : XOR2
      port map(A => AO6_70_Y, B => BUF_12_Y, Y => PP3_8_net);
    AOI1_E_1_inst : AOI1
      port map(A => XOR2_13_Y, B => OR3_2_Y, C => AND3_6_Y, Y => 
        E_1_net);
    XOR2_PP0_3_inst : XOR2
      port map(A => AO6_4_Y, B => BUF_26_Y, Y => PP0_3_net);
    AO6_66 : AO6
      port map(A => BUF_27_Y, B => AO16_13_Y, C => BUF_28_Y, D => 
        XOR2_25_Y, Y => AO6_66_Y);
    DF1_SumA_11_inst : DF1
      port map(D => FA1_72_CO, CLK => Clock, Q => SumA_11_net);
    DF1_62 : DF1
      port map(D => PP5_6_net, CLK => Clock, Q => DF1_62_Q);
    AO16_11 : AO16
      port map(A => DataB(5), B => DataB(6), C => BUF_12_Y, Y => 
        AO16_11_Y);
    XOR2_5 : XOR2
      port map(A => DataB(7), B => DataB(8), Y => XOR2_5_Y);
    HA1_4 : HA1
      port map(A => DF1_47_Q, B => VCC_1_net, CO => HA1_4_CO, 
        S => HA1_4_S);
    XOR2_PP4_6_inst : XOR2
      port map(A => AO6_89_Y, B => BUF_37_Y, Y => PP4_6_net);
    XOR2_PP0_8_inst : XOR2
      port map(A => AO6_38_Y, B => BUF_26_Y, Y => PP0_8_net);
    ADD1_Mult_29_inst : ADD1
      port map(A => SumA_28_net, B => SumB_28_net, FCI => 
        ADD1_Mult_28_FCO, S => Mult(29), FCO => ADD1_Mult_29_FCO);
    AO6_93 : AO6
      port map(A => BUF_1_Y, B => AO16_8_Y, C => BUF_32_Y, D => 
        XOR2_3_Y, Y => AO6_93_Y);
    FA1_59 : FA1
      port map(A => FA1_0_CO, B => FA1_13_S, CI => FA1_66_S, 
        CO => FA1_59_CO, S => FA1_59_S);
    ADD1_Mult_21_inst : ADD1
      port map(A => SumA_20_net, B => SumB_20_net, FCI => 
        ADD1_Mult_20_FCO, S => Mult(21), FCO => ADD1_Mult_21_FCO);
    AO6_21 : AO6
      port map(A => BUF_1_Y, B => AO16_6_Y, C => BUF_32_Y, D => 
        XOR2_18_Y, Y => AO6_21_Y);
    XOR2_PP0_7_inst : XOR2
      port map(A => AO6_63_Y, B => BUF_26_Y, Y => PP0_7_net);
    ADD1_Mult_15_inst : ADD1
      port map(A => SumA_14_net, B => SumB_14_net, FCI => 
        ADD1_Mult_14_FCO, S => Mult(15), FCO => ADD1_Mult_15_FCO);
    DF1_143 : DF1
      port map(D => PP0_4_net, CLK => Clock, Q => DF1_143_Q);
    AO6_92 : AO6
      port map(A => BUF_43_Y, B => AND2A_1_Y, C => BUF_42_Y, D => 
        DataB(0), Y => AO6_92_Y);
    FA1_71 : FA1
      port map(A => DF1_147_Q, B => DF1_45_Q, CI => DF1_46_Q, 
        CO => FA1_71_CO, S => FA1_71_S);
    FA1_93 : FA1
      port map(A => FA1_66_CO, B => FA1_33_S, CI => FA1_15_S, 
        CO => FA1_93_CO, S => FA1_93_S);
    XOR2_PP7_13_inst : XOR2
      port map(A => AO6_21_Y, B => BUF_20_Y, Y => PP7_13_net);
    AO6_109 : AO6
      port map(A => BUF_36_Y, B => AO16_12_Y, C => BUF_13_Y, D => 
        XOR2_2_Y, Y => AO6_109_Y);
    AO16_6 : AO16
      port map(A => DataB(13), B => DataB(14), C => BUF_20_Y, 
        Y => AO16_6_Y);
    BUF_1 : BUFF
      port map(A => DataA(12), Y => BUF_1_Y);
    FA1_77 : FA1
      port map(A => FA1_42_CO, B => HA1_6_S, CI => FA1_43_S, 
        CO => FA1_77_CO, S => FA1_77_S);
    BUF_2 : BUFF
      port map(A => DataA(4), Y => BUF_2_Y);
    XOR2_PP3_13_inst : XOR2
      port map(A => AO6_59_Y, B => BUF_3_Y, Y => PP3_13_net);
    MX2_3 : MX2
      port map(A => BUF_41_Y, B => XOR2_19_Y, S => XOR2_6_Y, Y => 
        MX2_3_Y);
    DF1_137 : DF1
      port map(D => PP0_13_net, CLK => Clock, Q => DF1_137_Q);
    ADD1_Mult_3_inst : ADD1
      port map(A => SumA_2_net, B => SumB_2_net, FCI => 
        ADD1_Mult_2_FCO, S => Mult(3), FCO => ADD1_Mult_3_FCO);
    XOR2_PP7_6_inst : XOR2
      port map(A => AO6_109_Y, B => BUF_22_Y, Y => PP7_6_net);
    AO6_31 : AO6
      port map(A => BUF_13_Y, B => AO16_12_Y, C => BUF_44_Y, D => 
        XOR2_2_Y, Y => AO6_31_Y);
    AO6_43 : AO6
      port map(A => BUF_28_Y, B => AO16_11_Y, C => BUF_39_Y, D => 
        XOR2_17_Y, Y => AO6_43_Y);
    DF1_71 : DF1
      port map(D => E_5_net, CLK => Clock, Q => DF1_71_Q);
    ADD1_Mult_1_inst : ADD1
      port map(A => SumA_0_net, B => SumB_0_net, FCI => 
        FCINIT_BUFF_0_FCO, S => Mult(1), FCO => ADD1_Mult_1_FCO);
    AO1_4 : AO1
      port map(A => XOR2_19_Y, B => OR3_3_Y, C => AND3_5_Y, Y => 
        AO1_4_Y);
    DF1_77 : DF1
      port map(D => PP2_3_net, CLK => Clock, Q => DF1_77_Q);
    DF1_107 : DF1
      port map(D => PP3_3_net, CLK => Clock, Q => DF1_107_Q);
    DF1_124 : DF1
      port map(D => PP0_5_net, CLK => Clock, Q => DF1_124_Q);
    AND2_2 : AND2
      port map(A => XOR2_25_Y, B => BUF_29_Y, Y => AND2_2_Y);
    AO6_10 : AO6
      port map(A => BUF_8_Y, B => AO16_1_Y, C => BUF_35_Y, D => 
        XOR2_10_Y, Y => AO6_10_Y);
    DF1_12 : DF1
      port map(D => PP6_14_net, CLK => Clock, Q => DF1_12_Q);
    ADD1_Mult_17_inst : ADD1
      port map(A => SumA_16_net, B => SumB_16_net, FCI => 
        ADD1_Mult_16_FCO, S => Mult(17), FCO => ADD1_Mult_17_FCO);
    XOR2_PP6_15_inst : XOR2
      port map(A => AO6_91_Y, B => BUF_6_Y, Y => PP6_15_net);
    AO6_42 : AO6
      port map(A => BUF_15_Y, B => AO16_2_Y, C => BUF_1_Y, D => 
        XOR2_6_Y, Y => AO6_42_Y);
    AND3_2 : AND3
      port map(A => DataB(3), B => DataB(4), C => DataB(5), Y => 
        AND3_2_Y);
    DF1_SumB_12_inst : DF1
      port map(D => FA1_73_S, CLK => Clock, Q => SumB_12_net);
    XOR2_PP7_7_inst : XOR2
      port map(A => AO6_31_Y, B => BUF_22_Y, Y => PP7_7_net);
    DF1_32 : DF1
      port map(D => PP6_15_net, CLK => Clock, Q => DF1_32_Q);
    DF1_130 : DF1
      port map(D => PP1_2_net, CLK => Clock, Q => DF1_130_Q);
    HA1_9 : HA1
      port map(A => DF1_93_Q, B => DF1_83_Q, CO => HA1_9_CO, S => 
        HA1_9_S);
    FA1_11 : FA1
      port map(A => FA1_85_CO, B => HA1_1_S, CI => FA1_67_S, 
        CO => FA1_11_CO, S => FA1_11_S);
    XOR2_12 : XOR2
      port map(A => AND2_7_Y, B => BUF_22_Y, Y => XOR2_12_Y);
    FA1_17 : FA1
      port map(A => FA1_36_CO, B => FA1_61_CO, CI => FA1_11_S, 
        CO => FA1_17_CO, S => FA1_17_S);
    AO16_2 : AO16
      port map(A => DataB(9), B => DataB(10), C => BUF_41_Y, Y => 
        AO16_2_Y);
    DF1_83 : DF1
      port map(D => PP6_5_net, CLK => Clock, Q => DF1_83_Q);
    DF1_100 : DF1
      port map(D => PP4_14_net, CLK => Clock, Q => DF1_100_Q);
    AO6_53 : AO6
      port map(A => BUF_1_Y, B => AO16_0_Y, C => BUF_32_Y, D => 
        XOR2_5_Y, Y => AO6_53_Y);
    OR3_7 : OR3
      port map(A => DataB(7), B => DataB(8), C => DataB(9), Y => 
        OR3_7_Y);
    AO6_118 : AO6
      port map(A => BUF_35_Y, B => AO16_12_Y, C => BUF_25_Y, D => 
        XOR2_2_Y, Y => AO6_118_Y);
    HA1_12 : HA1
      port map(A => DF1_152_Q, B => DF1_109_Q, CO => HA1_12_CO, 
        S => HA1_12_S);
    DF1_150 : DF1
      port map(D => PP5_3_net, CLK => Clock, Q => DF1_150_Q);
    BUF_37 : BUFF
      port map(A => DataB(9), Y => BUF_37_Y);
    AO6_15 : AO6
      port map(A => BUF_0_Y, B => AO16_7_Y, C => BUF_46_Y, D => 
        XOR2_28_Y, Y => AO6_15_Y);
    DF1_80 : DF1
      port map(D => PP7_4_net, CLK => Clock, Q => DF1_80_Q);
    XOR2_PP7_5_inst : XOR2
      port map(A => AO6_111_Y, B => BUF_22_Y, Y => PP7_5_net);
    XOR2_16 : XOR2
      port map(A => AND2_0_Y, B => BUF_26_Y, Y => XOR2_16_Y);
    FA1_41 : FA1
      port map(A => DF1_66_Q, B => DF1_15_Q, CI => DF1_121_Q, 
        CO => FA1_41_CO, S => FA1_41_S);
    FA1_96 : FA1
      port map(A => FA1_54_CO, B => FA1_37_S, CI => FA1_25_S, 
        CO => FA1_96_CO, S => FA1_96_S);
    DF1_135 : DF1
      port map(D => PP1_7_net, CLK => Clock, Q => DF1_135_Q);
    AO6_52 : AO6
      port map(A => BUF_25_Y, B => AO16_4_Y, C => BUF_4_Y, D => 
        XOR2_29_Y, Y => AO6_52_Y);
    XOR2_PP4_2_inst : XOR2
      port map(A => AO6_58_Y, B => BUF_37_Y, Y => PP4_2_net);
    DF1_SumB_21_inst : DF1
      port map(D => FA1_74_S, CLK => Clock, Q => SumB_21_net);
    XOR2_PP2_12_inst : XOR2
      port map(A => AO6_17_Y, B => BUF_30_Y, Y => PP2_12_net);
    DF1_85 : DF1
      port map(D => PP2_8_net, CLK => Clock, Q => DF1_85_Q);
    AO6_97 : AO6
      port map(A => BUF_8_Y, B => AO16_5_Y, C => BUF_35_Y, D => 
        XOR2_8_Y, Y => AO6_97_Y);
    FA1_81 : FA1
      port map(A => FA1_75_CO, B => HA1_7_S, CI => FA1_31_S, 
        CO => FA1_81_CO, S => FA1_81_S);
    FA1_47 : FA1
      port map(A => DF1_68_Q, B => DF1_75_Q, CI => DF1_56_Q, 
        CO => FA1_47_CO, S => FA1_47_S);
    FA1_94 : FA1
      port map(A => DF1_61_Q, B => DF1_140_Q, CI => DF1_85_Q, 
        CO => FA1_94_CO, S => FA1_94_S);
    DF1_2 : DF1
      port map(D => PP2_0_net, CLK => Clock, Q => DF1_2_Q);
    DF1_79 : DF1
      port map(D => PP1_5_net, CLK => Clock, Q => DF1_79_Q);
    FA1_87 : FA1
      port map(A => FA1_63_CO, B => DF1_1_Q, CI => FA1_71_S, 
        CO => FA1_87_CO, S => FA1_87_S);
    DF1_SumA_14_inst : DF1
      port map(D => FA1_96_CO, CLK => Clock, Q => SumA_14_net);
    DF1_105 : DF1
      port map(D => PP6_11_net, CLK => Clock, Q => DF1_105_Q);
    DF1_44 : DF1
      port map(D => PP5_9_net, CLK => Clock, Q => DF1_44_Q);
    DF1_52 : DF1
      port map(D => PP7_2_net, CLK => Clock, Q => DF1_52_Q);
    BUF_40 : BUFF
      port map(A => DataA(15), Y => BUF_40_Y);
    DF1_116 : DF1
      port map(D => E_7_net, CLK => Clock, Q => DF1_116_Q);
    AO6_98 : AO6
      port map(A => BUF_5_Y, B => AO16_13_Y, C => BUF_14_Y, D => 
        XOR2_25_Y, Y => AO6_98_Y);
    DF1_SumA_27_inst : DF1
      port map(D => FA1_91_CO, CLK => Clock, Q => SumA_27_net);
    FA1_58 : FA1
      port map(A => FA1_29_CO, B => HA1_15_CO, CI => FA1_14_S, 
        CO => FA1_58_CO, S => FA1_58_S);
    FA1_52 : FA1
      port map(A => HA1_14_CO, B => DF1_7_Q, CI => FA1_50_CO, 
        CO => FA1_52_CO, S => FA1_52_S);
    MX2_PP2_16_inst : MX2
      port map(A => MX2_0_Y, B => AO1_2_Y, S => AO16_9_Y, Y => 
        PP2_16_net);
    XOR2_PP0_10_inst : XOR2
      port map(A => AO6_48_Y, B => BUF_23_Y, Y => PP0_10_net);
    AO6_1 : AO6
      port map(A => BUF_14_Y, B => AO16_3_Y, C => BUF_10_Y, D => 
        XOR2_4_Y, Y => AO6_1_Y);
    AO6_113 : AO6
      port map(A => BUF_24_Y, B => AO16_3_Y, C => BUF_16_Y, D => 
        XOR2_4_Y, Y => AO6_113_Y);
    XOR2_PP6_2_inst : XOR2
      port map(A => AO6_64_Y, B => BUF_17_Y, Y => PP6_2_net);
    FA1_21 : FA1
      port map(A => DF1_35_Q, B => DF1_108_Q, CI => DF1_134_Q, 
        CO => FA1_21_CO, S => FA1_21_S);
    BUF_42 : BUFF
      port map(A => DataA(11), Y => BUF_42_Y);
    FA1_73 : FA1
      port map(A => FA1_7_CO, B => FA1_9_S, CI => FA1_54_S, CO => 
        FA1_73_CO, S => FA1_73_S);
    AND2_5 : AND2
      port map(A => XOR2_17_Y, B => BUF_29_Y, Y => AND2_5_Y);
    XOR2_28 : XOR2
      port map(A => DataB(5), B => DataB(6), Y => XOR2_28_Y);
    FA1_27 : FA1
      port map(A => FA1_67_CO, B => HA1_1_CO, CI => FA1_86_S, 
        CO => FA1_27_CO, S => FA1_27_S);
    XOR2_PP5_10_inst : XOR2
      port map(A => AO6_104_Y, B => BUF_41_Y, Y => PP5_10_net);
    DF1_SumB_10_inst : DF1
      port map(D => FA1_72_S, CLK => Clock, Q => SumB_10_net);
    AO6_47 : AO6
      port map(A => BUF_5_Y, B => AO16_10_Y, C => BUF_14_Y, D => 
        XOR2_21_Y, Y => AO6_47_Y);
    DF1_SumB_3_inst : DF1
      port map(D => FA1_84_S, CLK => Clock, Q => SumB_3_net);
    DF1_6 : DF1
      port map(D => PP4_1_net, CLK => Clock, Q => DF1_6_Q);
    XOR2_PP4_15_inst : XOR2
      port map(A => AO6_75_Y, B => BUF_33_Y, Y => PP4_15_net);
    XOR2_PP1_11_inst : XOR2
      port map(A => AO6_84_Y, B => BUF_11_Y, Y => PP1_11_net);
    BUF_9 : BUFF
      port map(A => DataA(10), Y => BUF_9_Y);
    XOR2_1 : XOR2
      port map(A => AND2_3_Y, B => BUF_17_Y, Y => XOR2_1_Y);
    DF1_SumB_15_inst : DF1
      port map(D => FA1_59_S, CLK => Clock, Q => SumB_15_net);
    XOR2_PP7_12_inst : XOR2
      port map(A => AO6_117_Y, B => BUF_20_Y, Y => PP7_12_net);
    AO6_48 : AO6
      port map(A => BUF_10_Y, B => AND2A_1_Y, C => BUF_43_Y, D => 
        DataB(0), Y => AO6_48_Y);
    XOR2_PP1_7_inst : XOR2
      port map(A => AO6_68_Y, B => BUF_18_Y, Y => PP1_7_net);
    BUF_17 : BUFF
      port map(A => DataB(13), Y => BUF_17_Y);
    XOR2_8 : XOR2
      port map(A => DataB(11), B => DataB(12), Y => XOR2_8_Y);
    BUF_27 : BUFF
      port map(A => DataA(2), Y => BUF_27_Y);
    XOR2_PP3_12_inst : XOR2
      port map(A => AO6_100_Y, B => BUF_3_Y, Y => PP3_12_net);
    FA1_31 : FA1
      port map(A => DF1_51_Q, B => DF1_77_Q, CI => DF1_142_Q, 
        CO => FA1_31_CO, S => FA1_31_S);
    ADD1_Mult_14_inst : ADD1
      port map(A => SumA_13_net, B => SumB_13_net, FCI => 
        ADD1_Mult_13_FCO, S => Mult(14), FCO => ADD1_Mult_14_FCO);
    DF1_48 : DF1
      port map(D => PP3_15_net, CLK => Clock, Q => DF1_48_Q);
    ADD1_Mult_2_inst : ADD1
      port map(A => SumA_1_net, B => SumB_1_net, FCI => 
        ADD1_Mult_1_FCO, S => Mult(2), FCO => ADD1_Mult_2_FCO);
    XOR2_PP5_5_inst : XOR2
      port map(A => AO6_50_Y, B => BUF_47_Y, Y => PP5_5_net);
    FA1_37 : FA1
      port map(A => HA1_0_CO, B => DF1_86_Q, CI => FA1_26_S, 
        CO => FA1_37_CO, S => FA1_37_S);
    XOR2_PP1_14_inst : XOR2
      port map(A => AO6_78_Y, B => BUF_11_Y, Y => PP1_14_net);
    AO6_57 : AO6
      port map(A => BUF_31_Y, B => AO16_2_Y, C => BUF_40_Y, D => 
        XOR2_6_Y, Y => AO6_57_Y);
    FA1_13 : FA1
      port map(A => FA1_24_CO, B => HA1_12_CO, CI => FA1_90_S, 
        CO => FA1_13_CO, S => FA1_13_S);
    ADD1_Mult_19_inst : ADD1
      port map(A => SumA_18_net, B => SumB_18_net, FCI => 
        ADD1_Mult_18_FCO, S => Mult(19), FCO => ADD1_Mult_19_FCO);
    AO6_14 : AO6
      port map(A => BUF_8_Y, B => AO16_12_Y, C => BUF_35_Y, D => 
        XOR2_2_Y, Y => AO6_14_Y);
    AO1_6 : AO1
      port map(A => XOR2_7_Y, B => OR3_0_Y, C => AND3_3_Y, Y => 
        AO1_6_Y);
    DF1_SumA_4_inst : DF1
      port map(D => FA1_84_CO, CLK => Clock, Q => SumA_4_net);
    XOR2_PP4_5_inst : XOR2
      port map(A => AO6_71_Y, B => BUF_37_Y, Y => PP4_5_net);
    XOR2_PP3_2_inst : XOR2
      port map(A => AO6_108_Y, B => BUF_12_Y, Y => PP3_2_net);
    ADD1_Mult_11_inst : ADD1
      port map(A => SumA_10_net, B => SumB_10_net, FCI => 
        ADD1_Mult_10_FCO, S => Mult(11), FCO => ADD1_Mult_11_FCO);
    DF1_92 : DF1
      port map(D => S_4_net, CLK => Clock, Q => DF1_92_Q);
    FA1_61 : FA1
      port map(A => FA1_41_CO, B => HA1_2_S, CI => FA1_85_S, 
        CO => FA1_61_CO, S => FA1_61_S);
    XOR2_PP5_7_inst : XOR2
      port map(A => AO6_28_Y, B => BUF_47_Y, Y => PP5_7_net);
    AND3_5 : AND3
      port map(A => DataB(9), B => DataB(10), C => DataB(11), 
        Y => AND3_5_Y);
    FA1_95 : FA1
      port map(A => FA1_25_CO, B => FA1_34_S, CI => FA1_0_S, 
        CO => FA1_95_CO, S => FA1_95_S);
    AO6_58 : AO6
      port map(A => BUF_35_Y, B => AO16_1_Y, C => BUF_25_Y, D => 
        XOR2_10_Y, Y => AO6_58_Y);
    DF1_121 : DF1
      port map(D => PP4_9_net, CLK => Clock, Q => DF1_121_Q);
    FA1_67 : FA1
      port map(A => DF1_76_Q, B => DF1_110_Q, CI => DF1_131_Q, 
        CO => FA1_67_CO, S => FA1_67_S);
    DF1_1 : DF1
      port map(D => PP7_0_net, CLK => Clock, Q => DF1_1_Q);
    AO6_70 : AO6
      port map(A => BUF_5_Y, B => AO16_11_Y, C => BUF_14_Y, D => 
        XOR2_17_Y, Y => AO6_70_Y);
    XOR2_PP7_2_inst : XOR2
      port map(A => AO6_118_Y, B => BUF_22_Y, Y => PP7_2_net);
    BUF_41 : BUFF
      port map(A => DataB(11), Y => BUF_41_Y);
    FA1_43 : FA1
      port map(A => DF1_115_Q, B => DF1_23_Q, CI => DF1_24_Q, 
        CO => FA1_43_CO, S => FA1_43_S);
    FA1_76 : FA1
      port map(A => FA1_57_CO, B => FA1_5_S, CI => FA1_7_S, CO => 
        FA1_76_CO, S => FA1_76_S);
    OR3_5 : OR3
      port map(A => DataB(5), B => DataB(6), C => DataB(7), Y => 
        OR3_5_Y);
    DF1_147 : DF1
      port map(D => PP2_10_net, CLK => Clock, Q => DF1_147_Q);
    XOR2_PP1_4_inst : XOR2
      port map(A => AO6_46_Y, B => BUF_18_Y, Y => PP1_4_net);
    AO6_19 : AO6
      port map(A => BUF_27_Y, B => AO16_10_Y, C => BUF_28_Y, D => 
        XOR2_21_Y, Y => AO6_19_Y);
    DF1_3 : DF1
      port map(D => PP6_1_net, CLK => Clock, Q => DF1_3_Q);
    DF1_128 : DF1
      port map(D => E_1_net, CLK => Clock, Q => DF1_128_Q);
    FA1_83 : FA1
      port map(A => DF1_13_Q, B => DF1_95_Q, CI => DF1_139_Q, 
        CO => FA1_83_CO, S => FA1_83_S);
    DF1_SumB_24_inst : DF1
      port map(D => FA1_69_S, CLK => Clock, Q => SumB_24_net);
    FA1_74 : FA1
      port map(A => FA1_48_CO, B => FA1_18_S, CI => FA1_92_S, 
        CO => FA1_74_CO, S => FA1_74_S);
    HA1_S_0_inst : HA1
      port map(A => XOR2_16_Y, B => DataB(1), CO => S_0_net, S => 
        PP0_0_net);
    AO6_80 : AO6
      port map(A => BUF_7_Y, B => AO16_10_Y, C => BUF_5_Y, D => 
        XOR2_21_Y, Y => AO6_80_Y);
    ADD1_Mult_31_inst : ADD1
      port map(A => SumA_30_net, B => SumB_30_net, FCI => 
        ADD1_Mult_30_FCO, S => Mult(31), FCO => ADD1_Mult_31_FCO);
    AND3_3 : AND3
      port map(A => DataB(11), B => DataB(12), C => DataB(13), 
        Y => AND3_3_Y);
    DF1_23 : DF1
      port map(D => PP0_16_net, CLK => Clock, Q => DF1_23_Q);
    AO6_91 : AO6
      port map(A => BUF_31_Y, B => AO16_8_Y, C => BUF_40_Y, D => 
        XOR2_3_Y, Y => AO6_91_Y);
    AO6_112 : AO6
      port map(A => BUF_25_Y, B => AO16_1_Y, C => BUF_4_Y, D => 
        XOR2_10_Y, Y => AO6_112_Y);
    AO16_10 : AO16
      port map(A => DataB(3), B => DataB(4), C => BUF_34_Y, Y => 
        AO16_10_Y);
    ADD1_Mult_8_inst : ADD1
      port map(A => SumA_7_net, B => SumB_7_net, FCI => 
        ADD1_Mult_7_FCO, S => Mult(8), FCO => ADD1_Mult_8_FCO);
    AO6_117 : AO6
      port map(A => BUF_15_Y, B => AO16_6_Y, C => BUF_1_Y, D => 
        XOR2_18_Y, Y => AO6_117_Y);
    AOI1_E_3_inst : AOI1
      port map(A => XOR2_15_Y, B => OR3_5_Y, C => AND3_4_Y, Y => 
        E_3_net);
    DF1_20 : DF1
      port map(D => PP1_8_net, CLK => Clock, Q => DF1_20_Q);
    AO6_75 : AO6
      port map(A => BUF_31_Y, B => AO16_0_Y, C => BUF_40_Y, D => 
        XOR2_5_Y, Y => AO6_75_Y);
    AO6_63 : AO6
      port map(A => BUF_7_Y, B => AND2A_0_Y, C => BUF_5_Y, D => 
        DataB(0), Y => AO6_63_Y);
    DF1_140 : DF1
      port map(D => PP0_12_net, CLK => Clock, Q => DF1_140_Q);
    FA1_23 : FA1
      port map(A => FA1_32_CO, B => FA1_28_S, CI => FA1_58_S, 
        CO => FA1_23_CO, S => FA1_23_S);
    MX2_PP4_16_inst : MX2
      port map(A => MX2_6_Y, B => AO1_0_Y, S => AO16_0_Y, Y => 
        PP4_16_net);
    ADD1_Mult_20_inst : ADD1
      port map(A => SumA_19_net, B => SumB_19_net, FCI => 
        ADD1_Mult_19_FCO, S => Mult(20), FCO => ADD1_Mult_20_FCO);
    DF1_122 : DF1
      port map(D => PP3_9_net, CLK => Clock, Q => DF1_122_Q);
    DF1_25 : DF1
      port map(D => PP0_2_net, CLK => Clock, Q => DF1_25_Q);
    AO1_5 : AO1
      port map(A => XOR2_13_Y, B => OR3_2_Y, C => AND3_6_Y, Y => 
        AO1_5_Y);
    DF1_SumB_19_inst : DF1
      port map(D => FA1_2_S, CLK => Clock, Q => SumB_19_net);
    DF1_113 : DF1
      port map(D => PP6_10_net, CLK => Clock, Q => DF1_113_Q);
    DF1_SumA_5_inst : DF1
      port map(D => FA1_82_CO, CLK => Clock, Q => SumA_5_net);
    DF1_84 : DF1
      port map(D => PP2_9_net, CLK => Clock, Q => DF1_84_Q);
    FA1_16 : FA1
      port map(A => FA1_92_CO, B => FA1_21_S, CI => FA1_45_S, 
        CO => FA1_16_CO, S => FA1_16_S);
    XOR2_PP2_3_inst : XOR2
      port map(A => AO6_19_Y, B => BUF_34_Y, Y => PP2_3_net);
    ADD1_Mult_26_inst : ADD1
      port map(A => SumA_25_net, B => SumB_25_net, FCI => 
        ADD1_Mult_25_FCO, S => Mult(26), FCO => ADD1_Mult_26_FCO);
    DF1_139 : DF1
      port map(D => PP5_7_net, CLK => Clock, Q => DF1_139_Q);
    AO6_85 : AO6
      port map(A => BUF_13_Y, B => AO16_1_Y, C => BUF_44_Y, D => 
        XOR2_10_Y, Y => AO6_85_Y);
    AOI1_E_5_inst : AOI1
      port map(A => XOR2_19_Y, B => OR3_3_Y, C => AND3_5_Y, Y => 
        E_5_net);
    AND3_6 : AND3
      port map(A => DataB(1), B => DataB(2), C => DataB(3), Y => 
        AND3_6_Y);
    MX2_5 : MX2
      port map(A => BUF_6_Y, B => XOR2_7_Y, S => XOR2_3_Y, Y => 
        MX2_5_Y);
    AO6_62 : AO6
      port map(A => BUF_39_Y, B => AO16_11_Y, C => BUF_45_Y, D => 
        XOR2_17_Y, Y => AO6_62_Y);
    DF1_5 : DF1
      port map(D => PP4_16_net, CLK => Clock, Q => DF1_5_Q);
    FA1_14 : FA1
      port map(A => DF1_144_Q, B => DF1_20_Q, CI => DF1_41_Q, 
        CO => FA1_14_CO, S => FA1_14_S);
    DF1_63 : DF1
      port map(D => PP0_11_net, CLK => Clock, Q => DF1_63_Q);
    AO6_41 : AO6
      port map(A => BUF_14_Y, B => AND2A_1_Y, C => BUF_10_Y, D => 
        DataB(0), Y => AO6_41_Y);
    AO6_20 : AO6
      port map(A => BUF_38_Y, B => AO16_0_Y, C => BUF_9_Y, D => 
        XOR2_5_Y, Y => AO6_20_Y);
    DF1_109 : DF1
      port map(D => PP6_3_net, CLK => Clock, Q => DF1_109_Q);
    BUF_35 : BUFF
      port map(A => DataA(1), Y => BUF_35_Y);
    DF1_46 : DF1
      port map(D => PP4_6_net, CLK => Clock, Q => DF1_46_Q);
end DEF_ARCH;
