------------------------------------------------------------------------------
--  This file is a part of the LPP VHDL IP LIBRARY
--  Copyright (C) 2009 - 2010, Laboratory of Plasmas Physic - CNRS
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
-------------------------------------------------------------------------------
--                    Author : Martin Morlot
--                   Mail : martin.morlot@lpp.polytechnique.fr
-------------------------------------------------------------------------------
library IEEE;
use IEEE.numeric_std.all;
use IEEE.std_logic_1164.all;

entity SelectInputs is
generic(
    Input_SZ : integer := 16);
port(
    clk     : in  std_logic;
    raz     : in  std_logic;
    Read    : in  std_logic;
    B1      : in std_logic_vector(Input_SZ-1 downto 0);
    B2      : in std_logic_vector(Input_SZ-1 downto 0);
    B3      : in std_logic_vector(Input_SZ-1 downto 0);
    E1      : in std_logic_vector(Input_SZ-1 downto 0);
    E2      : in std_logic_vector(Input_SZ-1 downto 0);
    Conjugate : out std_logic;
    Take    : out std_logic;
    ReadFIFO : out std_logic_vector(4 downto 0); --B1,B2,B3,E1,E2
    Statu : out std_logic_vector(3 downto 0);    
    OP1     : out std_logic_vector(Input_SZ-1 downto 0);    
    OP2     : out std_logic_vector(Input_SZ-1 downto 0)
);
end SelectInputs;


architecture ar_SelectInputs of SelectInputs is

signal Read_reg : std_logic;
signal i : integer range 0 to 128;
signal j : integer range 0 to 15;
signal Read_int : std_logic_vector(4 downto 0);

type state is (stX,sta,stb,st1,st2,idl1,idl2);
signal ect : state;

begin
    process(clk,raz)
    begin
    
        if(raz='0')then
            Take <= '0';
            i <= 0;
            j <= 0;
            Read_reg <= '0';
            ect <= stX;
        
        elsif(clk'event and clk='1')then
            Read_reg <= Read;
              
            case ect is

                when stX =>
                    i <= 1;                    
                    if(Read_reg='0' and Read='1')then
                        if(j=15)then
                            j <= 1;
                        else
                            j<= j+1;
                        end if;
                        ect <= idl1;
                    end if;                

                when idl1 =>
                    ect <= st1;                
                
                when st1 =>
                    Take <= '1';
                    ect <= sta;
                
                when sta =>                    
                    if(Read_reg='0' and Read='1')then
                        ect <= idl2;
                    end if;

                when idl2 =>
                    ect <= st2;
                
                when st2 =>
                    Take <= '0';
                    ect <= stb;
                
                when stb =>                    
                    if(i=128)then                        
                        ect <= stX;
                    elsif(Read_reg='0' and Read='1')then
                        i <= i+1;
                        ect <= idl1;                                            
                    end if;

            end case;
        end if;
    end process;

Statu <= std_logic_vector(to_unsigned(j,4));

with j select
    Read_int <= "10000" when 1,
                "11000" when 2,
                "01000" when 3,
                "10100" when 4,
                "01100" when 5,
                "00100" when 6,
                "10010" when 7,
                "01010" when 8,
                "00110" when 9,
                "00010" when 10,
                "10001" when 11,
                "01001" when 12,
                "00101" when 13,
                "00011" when 14,
                "00001" when 15,                
                "00000" when others;  

with ect select
    ReadFIFO <= Read_int when idl1,
                Read_int when idl2,
                "00000" when others;


with j select
    OP1 <=  B1 when 1,
            B1 when 2,
            B1 when 4,
            B1 when 7,
            B1 when 11,
            B2 when 3,
            B2 when 5,
            B2 when 8,
            B2 when 12,
            B3 when 6,
            B3 when 9,
            B3 when 13,
            E1 when 10,
            E1 when 14,
            E2 when 15,            
            X"FFFF" when others;


with j select
    OP2 <=  B1 when 1,
            B2 when 2,
            B2 when 3,
            B3 when 4,
            B3 when 5,
            B3 when 6,
            E1 when 7,
            E1 when 8,
            E1 when 9,
            E1 when 10,
            E2 when 11,
            E2 when 12,
            E2 when 13,
            E2 when 14,
            E2 when 15,
            X"FFFF" when others;


with j select 
    Conjugate <= '1' when 1,
                 '1' when 3,
                 '1' when 6,
                 '1' when 10,
                 '1' when 15,
                 '0' when others; 


end ar_SelectInputs;