--------------------------------------------------------------------------------
-- Copyright 2007 Actel Corporation.  All rights reserved.

-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
-- ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
-- IN ADVANCE IN WRITING.

-- Revision 3.0 April 30, 2007 : v3.0 CoreFFT Release
--  File:		twiddle.v
--
--  Description: CoreFFT
--               Twiddle factor table
--
--  Rev: 0.1 5/10/2005 8:36AM   VD  : Pre Production
--  History:		5/10/2005 8:36AM - created
--
--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE work.fft_components.all;

ENTITY twiddle IS
  PORT (
    A : IN std_logic_vector(gLOGPTS-2 DOWNTO 0);
    T : OUT std_logic_vector(gTDWIDTH-1 DOWNTO 0));
END ENTITY twiddle;

ARCHITECTURE translated OF twiddle IS
  SIGNAL T_int : std_logic_vector(gTDWIDTH-1 DOWNTO 0);

BEGIN
  T <= T_int;

  PROCESS (A)
    VARIABLE T_int1  : std_logic_vector(gTDWIDTH-1 DOWNTO 0);
  BEGIN
    CASE A IS      -- synopsys parallel_case
      WHEN "0000000" => T_int1 := "00000000000000000111111111111111"; -- X0000 X7fff
      WHEN "0000001" => T_int1 := "00000011001001000111111111110101"; -- X0324 X7ff5
      WHEN "0000010" => T_int1 := "00000110010010000111111111011000"; -- X0648 X7fd8
      WHEN "0000011" => T_int1 := "00001001011010100111111110100110"; -- X096a X7fa6
      WHEN "0000100" => T_int1 := "00001100100011000111111101100001"; -- X0c8c X7f61
      WHEN "0000101" => T_int1 := "00001111101010110111111100001001"; -- X0fab X7f09
      WHEN "0000110" => T_int1 := "00010010110010000111111010011100"; -- X12c8 X7e9c
      WHEN "0000111" => T_int1 := "00010101111000100111111000011101"; -- X15e2 X7e1d
      WHEN "0001000" => T_int1 := "00011000111110010111110110001001"; -- X18f9 X7d89
      WHEN "0001001" => T_int1 := "00011100000010110111110011100011"; -- X1c0b X7ce3
      WHEN "0001010" => T_int1 := "00011111000110100111110000101001"; -- X1f1a X7c29
      WHEN "0001011" => T_int1 := "00100010001000110111101101011100"; -- X2223 X7b5c
      WHEN "0001100" => T_int1 := "00100101001010000111101001111100"; -- X2528 X7a7c
      WHEN "0001101" => T_int1 := "00101000001001100111100110001001"; -- X2826 X7989
      WHEN "0001110" => T_int1 := "00101011000111110111100010000100"; -- X2b1f X7884
      WHEN "0001111" => T_int1 := "00101110000100010111011101101011"; -- X2e11 X776b
      WHEN "0010000" => T_int1 := "00110000111110110111011001000001"; -- X30fb X7641
      WHEN "0010001" => T_int1 := "00110011110111110111010100000100"; -- X33df X7504
      WHEN "0010010" => T_int1 := "00110110101110100111001110110101"; -- X36ba X73b5
      WHEN "0010011" => T_int1 := "00111001100011000111001001010100"; -- X398c X7254
      WHEN "0010100" => T_int1 := "00111100010101100111000011100010"; -- X3c56 X70e2
      WHEN "0010101" => T_int1 := "00111111000101110110111101011110"; -- X3f17 X6f5e
      WHEN "0010110" => T_int1 := "01000001110011100110110111001001"; -- X41ce X6dc9
      WHEN "0010111" => T_int1 := "01000100011110100110110000100011"; -- X447a X6c23
      WHEN "0011000" => T_int1 := "01000111000111000110101001101101"; -- X471c X6a6d
      WHEN "0011001" => T_int1 := "01001001101101000110100010100110"; -- X49b4 X68a6
      WHEN "0011010" => T_int1 := "01001100001111110110011011001111"; -- X4c3f X66cf
      WHEN "0011011" => T_int1 := "01001110101111110110010011101000"; -- X4ebf X64e8
      WHEN "0011100" => T_int1 := "01010001001100110110001011110001"; -- X5133 X62f1
      WHEN "0011101" => T_int1 := "01010011100110110110000011101011"; -- X539b X60eb
      WHEN "0011110" => T_int1 := "01010101111101010101111011010111"; -- X55f5 X5ed7
      WHEN "0011111" => T_int1 := "01011000010000100101110010110011"; -- X5842 X5cb3
      WHEN "0100000" => T_int1 := "01011010100000100101101010000010"; -- X5a82 X5a82
      WHEN "0100001" => T_int1 := "01011100101100110101100001000010"; -- X5cb3 X5842
      WHEN "0100010" => T_int1 := "01011110110101110101010111110101"; -- X5ed7 X55f5
      WHEN "0100011" => T_int1 := "01100000111010110101001110011011"; -- X60eb X539b
      WHEN "0100100" => T_int1 := "01100010111100010101000100110011"; -- X62f1 X5133
      WHEN "0100101" => T_int1 := "01100100111010000100111010111111"; -- X64e8 X4ebf
      WHEN "0100110" => T_int1 := "01100110110011110100110000111111"; -- X66cf X4c3f
      WHEN "0100111" => T_int1 := "01101000101001100100100110110100"; -- X68a6 X49b4
      WHEN "0101000" => T_int1 := "01101010011011010100011100011100"; -- X6a6d X471c
      WHEN "0101001" => T_int1 := "01101100001000110100010001111010"; -- X6c23 X447a
      WHEN "0101010" => T_int1 := "01101101110010010100000111001110"; -- X6dc9 X41ce
      WHEN "0101011" => T_int1 := "01101111010111100011111100010111"; -- X6f5e X3f17
      WHEN "0101100" => T_int1 := "01110000111000100011110001010110"; -- X70e2 X3c56
      WHEN "0101101" => T_int1 := "01110010010101000011100110001100"; -- X7254 X398c
      WHEN "0101110" => T_int1 := "01110011101101010011011010111010"; -- X73b5 X36ba
      WHEN "0101111" => T_int1 := "01110101000001000011001111011111"; -- X7504 X33df
      WHEN "0110000" => T_int1 := "01110110010000010011000011111011"; -- X7641 X30fb
      WHEN "0110001" => T_int1 := "01110111011010110010111000010001"; -- X776b X2e11
      WHEN "0110010" => T_int1 := "01111000100001000010101100011111"; -- X7884 X2b1f
      WHEN "0110011" => T_int1 := "01111001100010010010100000100110"; -- X7989 X2826
      WHEN "0110100" => T_int1 := "01111010011111000010010100101000"; -- X7a7c X2528
      WHEN "0110101" => T_int1 := "01111011010111000010001000100011"; -- X7b5c X2223
      WHEN "0110110" => T_int1 := "01111100001010010001111100011010"; -- X7c29 X1f1a
      WHEN "0110111" => T_int1 := "01111100111000110001110000001011"; -- X7ce3 X1c0b
      WHEN "0111000" => T_int1 := "01111101100010010001100011111001"; -- X7d89 X18f9
      WHEN "0111001" => T_int1 := "01111110000111010001010111100010"; -- X7e1d X15e2
      WHEN "0111010" => T_int1 := "01111110100111000001001011001000"; -- X7e9c X12c8
      WHEN "0111011" => T_int1 := "01111111000010010000111110101011"; -- X7f09 X0fab
      WHEN "0111100" => T_int1 := "01111111011000010000110010001100"; -- X7f61 X0c8c
      WHEN "0111101" => T_int1 := "01111111101001100000100101101010"; -- X7fa6 X096a
      WHEN "0111110" => T_int1 := "01111111110110000000011001001000"; -- X7fd8 X0648
      WHEN "0111111" => T_int1 := "01111111111101010000001100100100"; -- X7ff5 X0324
      WHEN "1000000" => T_int1 := "01111111111111110000000000000000"; -- X7fff X0000
      WHEN "1000001" => T_int1 := "01111111111101011111110011011100"; -- X7ff5 Xfcdc
      WHEN "1000010" => T_int1 := "01111111110110001111100110111000"; -- X7fd8 Xf9b8
      WHEN "1000011" => T_int1 := "01111111101001101111011010010110"; -- X7fa6 Xf696
      WHEN "1000100" => T_int1 := "01111111011000011111001101110100"; -- X7f61 Xf374
      WHEN "1000101" => T_int1 := "01111111000010011111000001010101"; -- X7f09 Xf055
      WHEN "1000110" => T_int1 := "01111110100111001110110100111000"; -- X7e9c Xed38
      WHEN "1000111" => T_int1 := "01111110000111011110101000011110"; -- X7e1d Xea1e
      WHEN "1001000" => T_int1 := "01111101100010011110011100000111"; -- X7d89 Xe707
      WHEN "1001001" => T_int1 := "01111100111000111110001111110101"; -- X7ce3 Xe3f5
      WHEN "1001010" => T_int1 := "01111100001010011110000011100110"; -- X7c29 Xe0e6
      WHEN "1001011" => T_int1 := "01111011010111001101110111011101"; -- X7b5c Xdddd
      WHEN "1001100" => T_int1 := "01111010011111001101101011011000"; -- X7a7c Xdad8
      WHEN "1001101" => T_int1 := "01111001100010011101011111011010"; -- X7989 Xd7da
      WHEN "1001110" => T_int1 := "01111000100001001101010011100001"; -- X7884 Xd4e1
      WHEN "1001111" => T_int1 := "01110111011010111101000111101111"; -- X776b Xd1ef
      WHEN "1010000" => T_int1 := "01110110010000011100111100000101"; -- X7641 Xcf05
      WHEN "1010001" => T_int1 := "01110101000001001100110000100001"; -- X7504 Xcc21
      WHEN "1010010" => T_int1 := "01110011101101011100100101000110"; -- X73b5 Xc946
      WHEN "1010011" => T_int1 := "01110010010101001100011001110100"; -- X7254 Xc674
      WHEN "1010100" => T_int1 := "01110000111000101100001110101010"; -- X70e2 Xc3aa
      WHEN "1010101" => T_int1 := "01101111010111101100000011101001"; -- X6f5e Xc0e9
      WHEN "1010110" => T_int1 := "01101101110010011011111000110010"; -- X6dc9 Xbe32
      WHEN "1010111" => T_int1 := "01101100001000111011101110000110"; -- X6c23 Xbb86
      WHEN "1011000" => T_int1 := "01101010011011011011100011100100"; -- X6a6d Xb8e4
      WHEN "1011001" => T_int1 := "01101000101001101011011001001100"; -- X68a6 Xb64c
      WHEN "1011010" => T_int1 := "01100110110011111011001111000001"; -- X66cf Xb3c1
      WHEN "1011011" => T_int1 := "01100100111010001011000101000001"; -- X64e8 Xb141
      WHEN "1011100" => T_int1 := "01100010111100011010111011001101"; -- X62f1 Xaecd
      WHEN "1011101" => T_int1 := "01100000111010111010110001100101"; -- X60eb Xac65
      WHEN "1011110" => T_int1 := "01011110110101111010101000001011"; -- X5ed7 Xaa0b
      WHEN "1011111" => T_int1 := "01011100101100111010011110111110"; -- X5cb3 Xa7be
      WHEN "1100000" => T_int1 := "01011010100000101010010101111110"; -- X5a82 Xa57e
      WHEN "1100001" => T_int1 := "01011000010000101010001101001101"; -- X5842 Xa34d
      WHEN "1100010" => T_int1 := "01010101111101011010000100101001"; -- X55f5 Xa129
      WHEN "1100011" => T_int1 := "01010011100110111001111100010101"; -- X539b X9f15
      WHEN "1100100" => T_int1 := "01010001001100111001110100001111"; -- X5133 X9d0f
      WHEN "1100101" => T_int1 := "01001110101111111001101100011000"; -- X4ebf X9b18
      WHEN "1100110" => T_int1 := "01001100001111111001100100110001"; -- X4c3f X9931
      WHEN "1100111" => T_int1 := "01001001101101001001011101011010"; -- X49b4 X975a
      WHEN "1101000" => T_int1 := "01000111000111001001010110010011"; -- X471c X9593
      WHEN "1101001" => T_int1 := "01000100011110101001001111011101"; -- X447a X93dd
      WHEN "1101010" => T_int1 := "01000001110011101001001000110111"; -- X41ce X9237
      WHEN "1101011" => T_int1 := "00111111000101111001000010100010"; -- X3f17 X90a2
      WHEN "1101100" => T_int1 := "00111100010101101000111100011110"; -- X3c56 X8f1e
      WHEN "1101101" => T_int1 := "00111001100011001000110110101100"; -- X398c X8dac
      WHEN "1101110" => T_int1 := "00110110101110101000110001001011"; -- X36ba X8c4b
      WHEN "1101111" => T_int1 := "00110011110111111000101011111100"; -- X33df X8afc
      WHEN "1110000" => T_int1 := "00110000111110111000100110111111"; -- X30fb X89bf
      WHEN "1110001" => T_int1 := "00101110000100011000100010010101"; -- X2e11 X8895
      WHEN "1110010" => T_int1 := "00101011000111111000011101111100"; -- X2b1f X877c
      WHEN "1110011" => T_int1 := "00101000001001101000011001110111"; -- X2826 X8677
      WHEN "1110100" => T_int1 := "00100101001010001000010110000100"; -- X2528 X8584
      WHEN "1110101" => T_int1 := "00100010001000111000010010100100"; -- X2223 X84a4
      WHEN "1110110" => T_int1 := "00011111000110101000001111010111"; -- X1f1a X83d7
      WHEN "1110111" => T_int1 := "00011100000010111000001100011101"; -- X1c0b X831d
      WHEN "1111000" => T_int1 := "00011000111110011000001001110111"; -- X18f9 X8277
      WHEN "1111001" => T_int1 := "00010101111000101000000111100011"; -- X15e2 X81e3
      WHEN "1111010" => T_int1 := "00010010110010001000000101100100"; -- X12c8 X8164
      WHEN "1111011" => T_int1 := "00001111101010111000000011110111"; -- X0fab X80f7
      WHEN "1111100" => T_int1 := "00001100100011001000000010011111"; -- X0c8c X809f
      WHEN "1111101" => T_int1 := "00001001011010101000000001011010"; -- X096a X805a
      WHEN "1111110" => T_int1 := "00000110010010001000000000101000"; -- X0648 X8028
      WHEN "1111111" => T_int1 := "00000011001001001000000000001011"; -- X0324 X800b
      WHEN OTHERS => NULL;
    END CASE;
    T_int <= T_int1;
  END PROCESS;

END ARCHITECTURE translated;
