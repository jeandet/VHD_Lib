



-----------------------------------------------------------------------------
-- LEON3 Demonstration design test bench configuration
-- Copyright (C) 2009 Aeroflex Gaisler
------------------------------------------------------------------------------


LIBRARY techmap;
USE techmap.gencomp.ALL;

PACKAGE config IS
-- Technology and synthesis options
  CONSTANT CFG_FABTECH        : INTEGER := inferred;
  CONSTANT CFG_MEMTECH        : INTEGER := inferred;
  --constant CFG_FABTECH : integer := apa3; --inferred;
  --constant CFG_MEMTECH : integer := apa3; --inferred;
  CONSTANT CFG_PADTECH        : INTEGER := inferred;
  CONSTANT CFG_NOASYNC        : INTEGER := 0;
  CONSTANT CFG_SCAN           : INTEGER := 0;
-- Clock generator
  CONSTANT CFG_CLKTECH        : INTEGER := inferred;
  CONSTANT CFG_CLKMUL         : INTEGER := 2;
  CONSTANT CFG_CLKDIV         : INTEGER := 2;
  CONSTANT CFG_OCLKDIV        : INTEGER := 1;
  CONSTANT CFG_OCLKBDIV       : INTEGER := 0;
  CONSTANT CFG_OCLKCDIV       : INTEGER := 0;
  CONSTANT CFG_PCIDLL         : INTEGER := 0;
  CONSTANT CFG_PCISYSCLK      : INTEGER := 0;
  CONSTANT CFG_CLK_NOFB       : INTEGER := 0;
-- LEON3 processor core
  CONSTANT CFG_LEON3          : INTEGER := 1;
  CONSTANT CFG_NCPU           : INTEGER := (1);
  CONSTANT CFG_NWIN           : INTEGER := (8);
  CONSTANT CFG_V8             : INTEGER := 0 + 4*0;
  CONSTANT CFG_MAC            : INTEGER := 0;
  CONSTANT CFG_BP             : INTEGER := 0;
  CONSTANT CFG_SVT            : INTEGER := 0;
  CONSTANT CFG_RSTADDR        : INTEGER := 16#00000#;
  CONSTANT CFG_LDDEL          : INTEGER := (1);
  CONSTANT CFG_NOTAG          : INTEGER := 0;
  CONSTANT CFG_NWP            : INTEGER := (0);
  CONSTANT CFG_PWD            : INTEGER := 0*2;
  CONSTANT CFG_FPU            : INTEGER := 0 + 16*0 + 32*0;
  CONSTANT CFG_GRFPUSH        : INTEGER := 0;
  CONSTANT CFG_ICEN           : INTEGER := 1;
  CONSTANT CFG_ISETS          : INTEGER := 1;
  CONSTANT CFG_ISETSZ         : INTEGER := 4;
  CONSTANT CFG_ILINE          : INTEGER := 8;
  CONSTANT CFG_IREPL          : INTEGER := 0;
  CONSTANT CFG_ILOCK          : INTEGER := 0;
  CONSTANT CFG_ILRAMEN        : INTEGER := 0;
  CONSTANT CFG_ILRAMADDR      : INTEGER := 16#8E#;
  CONSTANT CFG_ILRAMSZ        : INTEGER := 1;
  CONSTANT CFG_DCEN           : INTEGER := 1;
  CONSTANT CFG_DSETS          : INTEGER := 1;
  CONSTANT CFG_DSETSZ         : INTEGER := 4;
  CONSTANT CFG_DLINE          : INTEGER := 8;
  CONSTANT CFG_DREPL          : INTEGER := 0;
  CONSTANT CFG_DLOCK          : INTEGER := 0;
  CONSTANT CFG_DSNOOP         : INTEGER := 0 + 0 + 4*0;
  CONSTANT CFG_DFIXED         : INTEGER := 16#0#;
  CONSTANT CFG_DLRAMEN        : INTEGER := 0;
  CONSTANT CFG_DLRAMADDR      : INTEGER := 16#8F#;
  CONSTANT CFG_DLRAMSZ        : INTEGER := 1;
  CONSTANT CFG_MMUEN          : INTEGER := 1;
  CONSTANT CFG_ITLBNUM        : INTEGER := 8;
  CONSTANT CFG_DTLBNUM        : INTEGER := 8;
  CONSTANT CFG_TLB_TYPE       : INTEGER := 0 + 1*2;
  CONSTANT CFG_TLB_REP        : INTEGER := 1;
  CONSTANT CFG_MMU_PAGE       : INTEGER := 0;
  CONSTANT CFG_DSU            : INTEGER := 0;
  CONSTANT CFG_ITBSZ          : INTEGER := 0;
  CONSTANT CFG_ATBSZ          : INTEGER := 0;
  CONSTANT CFG_LEON3FT_EN     : INTEGER := 0;
  CONSTANT CFG_IUFT_EN        : INTEGER := 0;
  CONSTANT CFG_FPUFT_EN       : INTEGER := 0;
  CONSTANT CFG_RF_ERRINJ      : INTEGER := 0;
  CONSTANT CFG_CACHE_FT_EN    : INTEGER := 0;
  CONSTANT CFG_CACHE_ERRINJ   : INTEGER := 0;
  CONSTANT CFG_LEON3_NETLIST  : INTEGER := 0;
  CONSTANT CFG_DISAS          : INTEGER := 0 + 0;
  CONSTANT CFG_PCLOW          : INTEGER := 2;
-- AMBA settings
  CONSTANT CFG_DEFMST         : INTEGER := (0);
  CONSTANT CFG_RROBIN         : INTEGER := 1;
  CONSTANT CFG_SPLIT          : INTEGER := 0;
  CONSTANT CFG_FPNPEN         : INTEGER := 0;
  CONSTANT CFG_AHBIO          : INTEGER := 16#FFF#;
  CONSTANT CFG_APBADDR        : INTEGER := 16#800#;
  CONSTANT CFG_AHB_MON        : INTEGER := 0;
  CONSTANT CFG_AHB_MONERR     : INTEGER := 0;
  CONSTANT CFG_AHB_MONWAR     : INTEGER := 0;
  CONSTANT CFG_AHB_DTRACE     : INTEGER := 0;
-- DSU UART
  CONSTANT CFG_AHB_UART       : INTEGER := 1;
-- JTAG based DSU interface
  CONSTANT CFG_AHB_JTAG       : INTEGER := 0;
-- Ethernet DSU
  CONSTANT CFG_DSU_ETH        : INTEGER := 0 + 0 + 0;
  CONSTANT CFG_ETH_BUF        : INTEGER := 1;
  CONSTANT CFG_ETH_IPM        : INTEGER := 16#C0A8#;
  CONSTANT CFG_ETH_IPL        : INTEGER := 16#0033#;
  CONSTANT CFG_ETH_ENM        : INTEGER := 16#020000#;
  CONSTANT CFG_ETH_ENL        : INTEGER := 16#000009#;
-- PROM/SRAM controller
  CONSTANT CFG_SRCTRL         : INTEGER := 0;
  CONSTANT CFG_SRCTRL_PROMWS  : INTEGER := 0;
  CONSTANT CFG_SRCTRL_RAMWS   : INTEGER := 0;
  CONSTANT CFG_SRCTRL_IOWS    : INTEGER := 0;
  CONSTANT CFG_SRCTRL_RMW     : INTEGER := 0;
  CONSTANT CFG_SRCTRL_8BIT    : INTEGER := 0;
  CONSTANT CFG_SRCTRL_SRBANKS : INTEGER := 1;
  CONSTANT CFG_SRCTRL_BANKSZ  : INTEGER := 0;
  CONSTANT CFG_SRCTRL_ROMASEL : INTEGER := 0;
-- LEON2 memory controller
  CONSTANT CFG_MCTRL_LEON2    : INTEGER := 1;
  CONSTANT CFG_MCTRL_RAM8BIT  : INTEGER := 0;
  CONSTANT CFG_MCTRL_RAM16BIT : INTEGER := 0;
  CONSTANT CFG_MCTRL_5CS      : INTEGER := 0;
  CONSTANT CFG_MCTRL_SDEN     : INTEGER := 1;
  CONSTANT CFG_MCTRL_SEPBUS   : INTEGER := 0;
  CONSTANT CFG_MCTRL_INVCLK   : INTEGER := 0;
  CONSTANT CFG_MCTRL_SD64     : INTEGER := 0;
  CONSTANT CFG_MCTRL_PAGE     : INTEGER := 1 + 0;
-- SDRAM controller
  CONSTANT CFG_SDCTRL         : INTEGER := 0;
  CONSTANT CFG_SDCTRL_INVCLK  : INTEGER := 0;
  CONSTANT CFG_SDCTRL_SD64    : INTEGER := 0;
  CONSTANT CFG_SDCTRL_PAGE    : INTEGER := 0 + 0;
-- AHB ROM
  CONSTANT CFG_AHBROMEN       : INTEGER := 0;
  CONSTANT CFG_AHBROPIP       : INTEGER := 0;
  CONSTANT CFG_AHBRODDR       : INTEGER := 16#000#;
  CONSTANT CFG_ROMADDR        : INTEGER := 16#000#;
  CONSTANT CFG_ROMMASK        : INTEGER := 16#E00# + 16#000#;
-- AHB RAM
  CONSTANT CFG_AHBRAMEN       : INTEGER := 1;
  CONSTANT CFG_AHBRSZ         : INTEGER := 1;
  CONSTANT CFG_AHBRADDR       : INTEGER := 16#A00#;
-- Gaisler Ethernet core
  CONSTANT CFG_GRETH          : INTEGER := 0;
  CONSTANT CFG_GRETH1G        : INTEGER := 0;
  CONSTANT CFG_ETH_FIFO       : INTEGER := 8;

-- CAN 2.0 interface
  CONSTANT CFG_CAN         : INTEGER := 0;
  CONSTANT CFG_CANIO       : INTEGER := 16#0#;
  CONSTANT CFG_CANIRQ      : INTEGER := 0;
  CONSTANT CFG_CANLOOP     : INTEGER := 0;
  CONSTANT CFG_CAN_SYNCRST : INTEGER := 0;
  CONSTANT CFG_CANFT       : INTEGER := 0;

-- PCI interface
  CONSTANT CFG_PCI      : INTEGER := 0;
  CONSTANT CFG_PCIVID   : INTEGER := 16#0#;
  CONSTANT CFG_PCIDID   : INTEGER := 16#0#;
  CONSTANT CFG_PCIDEPTH : INTEGER := 8;
  CONSTANT CFG_PCI_MTF  : INTEGER := 1;

-- PCI arbiter
  CONSTANT CFG_PCI_ARB      : INTEGER := 0;
  CONSTANT CFG_PCI_ARBAPB   : INTEGER := 0;
  CONSTANT CFG_PCI_ARB_NGNT : INTEGER := 4;

-- PCI trace buffer
  CONSTANT CFG_PCITBUFEN : INTEGER := 0;
  CONSTANT CFG_PCITBUF   : INTEGER := 256;

-- Spacewire interface
  CONSTANT CFG_SPW_EN       : INTEGER := 0;
  CONSTANT CFG_SPW_NUM      : INTEGER := 1;
  CONSTANT CFG_SPW_AHBFIFO  : INTEGER := 4;
  CONSTANT CFG_SPW_RXFIFO   : INTEGER := 16;
  CONSTANT CFG_SPW_RMAP     : INTEGER := 0;
  CONSTANT CFG_SPW_RMAPBUF  : INTEGER := 4;
  CONSTANT CFG_SPW_RMAPCRC  : INTEGER := 0;
  CONSTANT CFG_SPW_NETLIST  : INTEGER := 0;
  CONSTANT CFG_SPW_FT       : INTEGER := 0;
  CONSTANT CFG_SPW_GRSPW    : INTEGER := 2;
  CONSTANT CFG_SPW_RXUNAL   : INTEGER := 0;
  CONSTANT CFG_SPW_DMACHAN  : INTEGER := 1;
  CONSTANT CFG_SPW_PORTS    : INTEGER := 1;
  CONSTANT CFG_SPW_INPUT    : INTEGER := 2;
  CONSTANT CFG_SPW_OUTPUT   : INTEGER := 0;
  CONSTANT CFG_SPW_RTSAME   : INTEGER := 0;
-- UART 1
  CONSTANT CFG_UART1_ENABLE : INTEGER := 1;
  CONSTANT CFG_UART1_FIFO   : INTEGER := 4;

-- UART 2
  CONSTANT CFG_UART2_ENABLE : INTEGER := 0;
  CONSTANT CFG_UART2_FIFO   : INTEGER := 1;

-- LEON3 interrupt controller
  CONSTANT CFG_IRQ3_ENABLE : INTEGER := 1;
  CONSTANT CFG_IRQ3_NSEC   : INTEGER := 0;

-- Modular timer
  CONSTANT CFG_GPT_ENABLE : INTEGER := 1;
  CONSTANT CFG_GPT_NTIM   : INTEGER := (2);
  CONSTANT CFG_GPT_SW     : INTEGER := (8);
  CONSTANT CFG_GPT_TW     : INTEGER := (32);
  CONSTANT CFG_GPT_IRQ    : INTEGER := (8);
  CONSTANT CFG_GPT_SEPIRQ : INTEGER := 1;
  CONSTANT CFG_GPT_WDOGEN : INTEGER := 1;
  CONSTANT CFG_GPT_WDOG   : INTEGER := 16#FFFF#;

-- GPIO port
  CONSTANT CFG_GRGPIO_ENABLE : INTEGER := 1;
  CONSTANT CFG_GRGPIO_IMASK  : INTEGER := 16#0000#;
  CONSTANT CFG_GRGPIO_WIDTH  : INTEGER := (8);

-- GRLIB debugging
  CONSTANT CFG_DUART : INTEGER := 1;
END;
