-- Version: 9.1 SP5 9.1.5.1

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_top_apbreg is

    port( status_full_ack    : out   std_logic_vector(3 downto 0);
          prdata_c           : out   std_logic_vector(31 downto 0);
          pirq_c             : out   std_logic_vector(15 to 15);
          addr_data_f2       : out   std_logic_vector(31 downto 0);
          status_new_err_3   : in    std_logic;
          status_new_err_0_2 : in    std_logic;
          status_new_err_0_0 : in    std_logic;
          status_new_err_0_1 : in    std_logic;
          status_full_err_0  : in    std_logic_vector(3 downto 0);
          status_full        : in    std_logic_vector(3 downto 0);
          addr_data_f3       : out   std_logic_vector(31 downto 0);
          nb_burst_available : out   std_logic_vector(10 downto 0);
          addr_data_f1       : out   std_logic_vector(31 downto 0);
          delta_f2_f1        : out   std_logic_vector(9 downto 0);
          addr_data_f0       : out   std_logic_vector(31 downto 0);
          delta_f2_f0        : out   std_logic_vector(9 downto 0);
          delta_snapshot     : out   std_logic_vector(15 downto 0);
          nb_snapshot_param  : out   std_logic_vector(10 downto 0);
          apbi_c_81          : in    std_logic;
          apbi_c_80          : in    std_logic;
          apbi_c_79          : in    std_logic;
          apbi_c_78          : in    std_logic;
          apbi_c_77          : in    std_logic;
          apbi_c_76          : in    std_logic;
          apbi_c_75          : in    std_logic;
          apbi_c_74          : in    std_logic;
          apbi_c_73          : in    std_logic;
          apbi_c_72          : in    std_logic;
          apbi_c_71          : in    std_logic;
          apbi_c_70          : in    std_logic;
          apbi_c_69          : in    std_logic;
          apbi_c_68          : in    std_logic;
          apbi_c_67          : in    std_logic;
          apbi_c_66          : in    std_logic;
          apbi_c_65          : in    std_logic;
          apbi_c_64          : in    std_logic;
          apbi_c_63          : in    std_logic;
          apbi_c_62          : in    std_logic;
          apbi_c_61          : in    std_logic;
          apbi_c_60          : in    std_logic;
          apbi_c_59          : in    std_logic;
          apbi_c_58          : in    std_logic;
          apbi_c_57          : in    std_logic;
          apbi_c_56          : in    std_logic;
          apbi_c_55          : in    std_logic;
          apbi_c_24          : in    std_logic;
          apbi_c_23          : in    std_logic;
          apbi_c_0           : in    std_logic;
          apbi_c_50          : in    std_logic;
          apbi_c_51          : in    std_logic;
          apbi_c_52          : in    std_logic;
          apbi_c_16          : in    std_logic;
          apbi_c_49          : in    std_logic;
          apbi_c_22          : in    std_logic;
          apbi_c_20          : in    std_logic;
          apbi_c_19          : in    std_logic;
          apbi_c_21          : in    std_logic;
          apbi_c_54          : in    std_logic;
          apbi_c_53          : in    std_logic;
          data_shaping_R0    : out   std_logic;
          data_shaping_R1    : out   std_logic;
          enable_f0          : out   std_logic;
          data_shaping_BW_c  : out   std_logic;
          burst_f2           : out   std_logic;
          burst_f1           : out   std_logic;
          burst_f0           : out   std_logic;
          enable_f3          : out   std_logic;
          enable_f2          : out   std_logic;
          data_shaping_SP1   : out   std_logic;
          enable_f1          : out   std_logic;
          data_shaping_SP0   : out   std_logic;
          data_shaping_R1_0  : out   std_logic;
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic;
          data_shaping_R0_0  : out   std_logic
        );

end lpp_top_apbreg;

architecture DEF_ARCH of lpp_top_apbreg is 

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal data_shaping_BW_1_sqmuxa, prdata_9_sqmuxa_0, N_931, 
        prdata_10_sqmuxa_0, prdata_12_sqmuxa_0, N_168, N_157, 
        N_933_0, N_930, addr_matrix_f0_0_1_sqmuxa_0, N_159, N_928, 
        addr_matrix_f0_1_1_sqmuxa_0, N_166, 
        addr_matrix_f1_1_sqmuxa_0, N_172, 
        addr_matrix_f2_1_sqmuxa_0, un1_apbi_2, 
        addr_data_f0_1_sqmuxa_0, addr_data_f1_1_sqmuxa_0, 
        addr_data_f2_1_sqmuxa_0, addr_data_f3_1_sqmuxa_0, N_161_0, 
        prdata_2_sqmuxa_0, prdata_3_sqmuxa_0, prdata_4_sqmuxa_0, 
        prdata_5_sqmuxa_0, N_168_0, \prdata_39_0_iv_14[4]\, 
        \nb_burst_available_m_i[4]\, \prdata_39_0_iv_9[4]\, 
        data_shaping_R1_m_i, \prdata_39_0_iv_11[4]\, 
        \prdata_39_0_iv_3[4]\, burst_f0_m_i, 
        \prdata_39_0_iv_7[4]\, \prdata_39_0_iv_10[4]\, 
        prdata_18_sqmuxa, \prdata_39_0_iv_6[4]\, 
        \addr_data_f3_m_i[4]\, \addr_data_f2_m_i[4]\, 
        \prdata_39_0_iv_5[4]\, prdata_14_sqmuxa, 
        \prdata_39_0_iv_2[4]\, \addr_matrix_f0_1_m_i[4]\, 
        \addr_matrix_f0_0_m_i[4]\, \prdata_39_0_iv_1[4]\, 
        prdata_16_sqmuxa, \delta_f2_f1_m_i[4]\, 
        \addr_data_f1_m_i[4]\, \status_full_err[0]\, 
        prdata_13_sqmuxa, 
        status_error_anticipating_empty_fifo_m_i, 
        \addr_matrix_f1[4]\, \addr_matrix_f2_m_i[4]\, 
        \prdata_39_0_iv_13[3]\, \nb_snapshot_param_m_i[3]\, 
        \prdata_39_0_iv_6[3]\, \prdata_39_0_iv_11[3]\, 
        \prdata_39_0_iv_12[3]\, \prdata_39_0_iv_3[3]\, 
        \prdata_39_0_iv_2[3]\, \prdata_39_0_iv_9[3]\, 
        \delta_snapshot_m_i[3]\, \prdata_39_0_iv_1[3]\, 
        \nb_burst_available_m_i[3]\, \delta_f2_f0_m_i[3]\, 
        \addr_data_f3_m_i[3]\, \prdata_39_0_iv_5[3]\, 
        \addr_matrix_f0_1_m_i[3]\, \addr_matrix_f0_0_m_i[3]\, 
        \status_full_m_i[3]\, prdata_15_sqmuxa, enable_f3_m_i, 
        \addr_data_f2_m_i[3]\, status_ready_matrix_f2_m_i, 
        \addr_matrix_f1[3]\, \addr_matrix_f2_m_i[3]\, 
        \prdata_39_0_iv_14[1]\, \prdata_39_0_iv_7[1]\, 
        \prdata_39_0_iv_6[1]\, \prdata_39_0_iv_10[1]\, 
        \prdata_39_0_iv_13[1]\, \prdata_39_0_iv_4[1]\, 
        \prdata_39_0_iv_3[1]\, data_shaping_SP0_m_i, 
        \prdata_39_0_iv_12[1]\, prdata_17_sqmuxa, 
        \prdata_39_0_iv_8[1]\, \prdata_39_0_iv_5[1]\, 
        enable_f1_m_i, \addr_matrix_f2_m_i[1]\, 
        \addr_matrix_f1_m_i[1]\, \prdata_39_0_iv_2[1]\, 
        \addr_matrix_f0_1_m_i[1]\, \addr_matrix_f0_0_m_i[1]\, 
        \status_full_m_i[1]\, \delta_f2_f1_m_i[1]\, 
        \addr_data_f2_m_i[1]\, \addr_data_f1_m_i[1]\, 
        prdata_0_sqmuxa, config_active_interruption_onError, 
        status_ready_matrix_f0_1_m_i, \prdata_39_0_iv_13[2]\, 
        \prdata_39_0_iv_6[2]\, \nb_snapshot_param_m_i[2]\, 
        data_shaping_SP1_m_i, \prdata_39_0_iv_12[2]\, 
        \prdata_39_0_iv_3[2]\, \prdata_39_0_iv_2[2]\, 
        \prdata_39_0_iv_9[2]\, \prdata_39_0_iv_11[2]\, 
        \prdata_39_0_iv_7[2]\, \status_full_m_i[2]\, 
        \delta_f2_f1_m_i[2]\, \prdata_39_0_iv_4[2]\, 
        enable_f2_m_i, \addr_matrix_f0_1_m_i[2]\, 
        \addr_matrix_f0_0_m_i[2]\, \prdata_39_0_iv_1[2]\, 
        \delta_f2_f0_m_i[2]\, \addr_data_f2_m_i[2]\, 
        status_ready_matrix_f1_m_i, \addr_matrix_f1[2]\, 
        \addr_matrix_f2_m_i[2]\, \prdata_39_0_iv_12[5]\, 
        \prdata_39_0_iv_5[5]\, \prdata_39_0_iv_4[5]\, 
        \nb_burst_available_m_i[5]\, \prdata_39_0_iv_11[5]\, 
        \prdata_39_0_iv_3[5]\, burst_f1_m_i, 
        \prdata_39_0_iv_7[5]\, \prdata_39_0_iv_10[5]\, 
        \prdata_39_0_iv_6[5]\, \prdata_39_0_iv_2[5]\, 
        \addr_matrix_f0_1_m_i[5]\, \addr_matrix_f0_0_m_i[5]\, 
        \prdata_39_0_iv_1[5]\, \delta_f2_f1_m_i[5]\, 
        \addr_data_f2_m_i[5]\, \addr_data_f1_m_i[5]\, 
        \status_full_err[1]\, 
        status_error_bad_component_error_m_i, \addr_matrix_f1[5]\, 
        \addr_matrix_f2_m_i[5]\, \prdata_39_0_iv_10[8]\, 
        \prdata_39_0_iv_3[8]\, \prdata_39_0_iv_2[8]\, 
        \nb_burst_available_m_i[8]\, \prdata_39_0_iv_9[8]\, 
        \prdata_39_0_iv_0[8]\, \delta_f2_f1_m_i[8]\, 
        \prdata_39_0_iv_6[8]\, \prdata_39_0_iv_8[8]\, 
        \delta_f2_f0_m_i[8]\, \addr_data_f3_m_i[8]\, 
        \nb_snapshot_param_m_i[8]\, \addr_matrix_f2_m_i[8]\, 
        \addr_matrix_f1_m_i[8]\, \delta_snapshot_m_i[8]\, 
        \addr_data_f2_m_i[8]\, \status_new_err[0]\, 
        \addr_data_f0_m_i[8]\, \addr_matrix_f0_0[8]\, 
        \addr_matrix_f0_1_m_i[8]\, \prdata_39_0_iv_14[0]\, 
        \prdata_39_0_iv_4[0]\, \prdata_39_0_iv_3[0]\, 
        \prdata_39_0_iv_11[0]\, \prdata_39_0_iv_13[0]\, 
        \delta_snapshot_m_i[0]\, \prdata_39_0_iv_2[0]\, 
        \prdata_39_0_iv_9[0]\, \prdata_39_0_iv_12[0]\, 
        \prdata_39_0_iv_7[0]\, \status_full_m_i[0]\, 
        \delta_f2_f1_m_i[0]\, \prdata_39_0_iv_5[0]\, 
        enable_f0_m_i, \addr_matrix_f0_1_m_i[0]\, 
        \addr_matrix_f0_0_m_i[0]\, \prdata_39_0_iv_1[0]\, 
        data_shaping_BW_m_i, \addr_data_f2_m_i[0]\, 
        \addr_data_f1_m_i[0]\, 
        config_active_interruption_onNewMatrix, 
        status_ready_matrix_f0_0_m_i, \addr_matrix_f1[0]\, 
        \addr_matrix_f2_m_i[0]\, \prdata_39_0_iv_11[6]\, 
        \prdata_39_0_iv_3[6]\, \prdata_39_0_iv_2[6]\, 
        \prdata_39_0_iv_8[6]\, \prdata_39_0_iv_10[6]\, 
        \prdata_39_0_iv_6[6]\, \prdata_39_0_iv_9[6]\, 
        \prdata_39_0_iv_5[6]\, \delta_f2_f0_m_i[6]\, 
        \addr_data_f3_m_i[6]\, burst_f2_m_i, 
        \addr_matrix_f2_m_i[6]\, \addr_matrix_f1_m_i[6]\, 
        \delta_snapshot_m_i[6]\, \addr_matrix_f0_1_m_i[6]\, 
        \addr_matrix_f0_0_m_i[6]\, \delta_f2_f1_m_i[6]\, 
        \addr_data_f2_m_i[6]\, \status_full_err[2]\, 
        \addr_data_f0_m_i[6]\, \prdata_39_0_iv_10[7]\, 
        \prdata_39_0_iv_3[7]\, \prdata_39_0_iv_2[7]\, 
        \nb_burst_available_m_i[7]\, \prdata_39_0_iv_9[7]\, 
        \delta_snapshot_m_i[7]\, \prdata_39_0_iv_1[7]\, 
        \prdata_39_0_iv_5[7]\, \prdata_39_0_iv_8[7]\, 
        \delta_f2_f0_m_i[7]\, \addr_data_f3_m_i[7]\, 
        \nb_snapshot_param_m_i[7]\, \addr_matrix_f0_1_m_i[7]\, 
        \addr_matrix_f0_0_m_i[7]\, \delta_f2_f1_m_i[7]\, 
        \addr_data_f2_m_i[7]\, \status_full_err[3]\, 
        \addr_data_f0_m_i[7]\, \addr_matrix_f1[7]\, 
        \addr_matrix_f2_m_i[7]\, \prdata_39_0_iv_10[9]\, 
        \prdata_39_0_iv_3[9]\, \prdata_39_0_iv_2[9]\, 
        \nb_burst_available_m_i[9]\, \prdata_39_0_iv_9[9]\, 
        \delta_snapshot_m_i[9]\, \prdata_39_0_iv_1[9]\, 
        \prdata_39_0_iv_5[9]\, \prdata_39_0_iv_8[9]\, 
        \delta_f2_f0_m_i[9]\, \addr_data_f3_m_i[9]\, 
        \nb_snapshot_param_m_i[9]\, \addr_matrix_f0_1_m_i[9]\, 
        \addr_matrix_f0_0_m_i[9]\, \delta_f2_f1_m_i[9]\, 
        \addr_data_f2_m_i[9]\, \status_new_err[1]\, 
        \addr_data_f0_m_i[9]\, \addr_matrix_f1[9]\, 
        \addr_matrix_f2_m_i[9]\, \prdata_39_0_iv_8[10]\, 
        \prdata_39_0_iv_2[10]\, \nb_snapshot_param_m_i[10]\, 
        \prdata_39_0_iv_5[10]\, \prdata_39_0_iv_7[10]\, 
        \prdata_39_0_iv_0[10]\, \addr_data_f3_m_i[10]\, 
        \prdata_39_0_iv_3[10]\, \prdata_39_0_iv_1[10]\, 
        \addr_data_f2_m_i[10]\, \status_new_err[2]\, 
        \addr_data_f0_m_i[10]\, \addr_matrix_f1[10]\, 
        \addr_matrix_f2_m_i[10]\, \addr_matrix_f0_0[10]\, 
        \addr_matrix_f0_1_m_i[10]\, \prdata_39_0_iv_6[11]\, 
        \addr_data_f0_m_i[11]\, \status_new_err_m_i[3]\, 
        \prdata_39_0_iv_3[11]\, \prdata_39_0_iv_5[11]\, 
        \prdata_39_0_iv_1[11]\, \prdata_39_0_iv_4[11]\, 
        \addr_matrix_f0_1_m_i[11]\, \addr_matrix_f0_0_m_i[11]\, 
        \addr_data_f3_m_i[11]\, \addr_data_f2_m_i[11]\, 
        \addr_matrix_f1[11]\, \addr_matrix_f2_m_i[11]\, 
        \prdata_39_0_iv_6[12]\, \prdata_39_0_iv_1[12]\, 
        \prdata_39_0_iv_0[12]\, \prdata_39_0_iv_3[12]\, 
        \addr_data_f2_m_i[12]\, \prdata_39_0_iv_2[12]\, 
        \addr_data_f1_m_i[12]\, \addr_matrix_f1[12]\, 
        \addr_matrix_f2_m_i[12]\, \addr_matrix_f0_0[12]\, 
        \addr_matrix_f0_1_m_i[12]\, \prdata_39_0_iv_6[13]\, 
        \prdata_39_0_iv_1[13]\, \prdata_39_0_iv_0[13]\, 
        \prdata_39_0_iv_3[13]\, \addr_data_f2_m_i[13]\, 
        \prdata_39_0_iv_2[13]\, \addr_data_f1_m_i[13]\, 
        \addr_matrix_f1[13]\, \addr_matrix_f2_m_i[13]\, 
        \addr_matrix_f0_0[13]\, \addr_matrix_f0_1_m_i[13]\, 
        \prdata_39_0_iv_6[14]\, \prdata_39_0_iv_1[14]\, 
        \prdata_39_0_iv_0[14]\, \prdata_39_0_iv_3[14]\, 
        \addr_data_f2_m_i[14]\, \prdata_39_0_iv_2[14]\, 
        \addr_data_f1_m_i[14]\, \addr_matrix_f1[14]\, 
        \addr_matrix_f2_m_i[14]\, \addr_matrix_f0_0[14]\, 
        \addr_matrix_f0_1_m_i[14]\, \prdata_39_0_iv_5[15]\, 
        \addr_data_f1_m_i[15]\, \addr_data_f0_m_i[15]\, 
        \delta_snapshot_m_i[15]\, \prdata_39_0_iv_4[15]\, 
        \addr_matrix_f0_1_m_i[15]\, \addr_matrix_f0_0_m_i[15]\, 
        \prdata_39_0_iv_1[15]\, \prdata_39_0_iv_3[15]\, 
        \addr_data_f2_m_i[15]\, \addr_matrix_f1[15]\, 
        \addr_matrix_f2_m_i[15]\, \prdata_39_0_iv_4[16]\, 
        \addr_matrix_f0_1_m_i[16]\, \addr_matrix_f0_0_m_i[16]\, 
        \prdata_39_0_iv_1[16]\, \prdata_39_0_iv_3[16]\, 
        \addr_data_f2_m_i[16]\, \prdata_39_0_iv_2[16]\, 
        \addr_data_f1_m_i[16]\, \addr_matrix_f1[16]\, 
        \addr_matrix_f2_m_i[16]\, \prdata_39_0_iv_4[17]\, 
        \addr_matrix_f0_1_m_i[17]\, \addr_matrix_f0_0_m_i[17]\, 
        \prdata_39_0_iv_1[17]\, \prdata_39_0_iv_3[17]\, 
        \addr_data_f2_m_i[17]\, \prdata_39_0_iv_2[17]\, 
        \addr_data_f1_m_i[17]\, \addr_matrix_f1[17]\, 
        \addr_matrix_f2_m_i[17]\, \prdata_39_0_iv_5[18]\, 
        \addr_data_f3_m_i[18]\, \addr_data_f2_m_i[18]\, 
        \prdata_39_0_iv_2[18]\, \addr_data_f1_m_i[18]\, 
        \prdata_39_0_iv_1[18]\, \addr_matrix_f1[18]\, 
        \addr_matrix_f2_m_i[18]\, \prdata_39_0_iv_0[18]\, 
        \addr_matrix_f0_0[18]\, \addr_matrix_f0_1_m_i[18]\, 
        \prdata_39_0_iv_4[19]\, \addr_matrix_f0_1_m_i[19]\, 
        \addr_matrix_f0_0_m_i[19]\, \prdata_39_0_iv_1[19]\, 
        \prdata_39_0_iv_3[19]\, \addr_data_f2_m_i[19]\, 
        \prdata_39_0_iv_2[19]\, \addr_data_f1_m_i[19]\, 
        prdata_4_sqmuxa, \addr_matrix_f1[19]\, 
        \addr_matrix_f2_m_i[19]\, \prdata_39_0_iv_4[20]\, 
        \addr_matrix_f0_1_m_i[20]\, \addr_matrix_f0_0_m_i[20]\, 
        \prdata_39_0_iv_1[20]\, \prdata_39_0_iv_3[20]\, 
        \addr_data_f2_m_i[20]\, \prdata_39_0_iv_2[20]\, 
        \addr_data_f1_m_i[20]\, \addr_matrix_f1[20]\, 
        \addr_matrix_f2_m_i[20]\, \prdata_39_0_iv_5[21]\, 
        \addr_data_f3_m_i[21]\, \addr_data_f2_m_i[21]\, 
        \prdata_39_0_iv_2[21]\, \addr_data_f1_m_i[21]\, 
        \prdata_39_0_iv_1[21]\, \addr_matrix_f1[21]\, 
        \addr_matrix_f2_m_i[21]\, \prdata_39_0_iv_0[21]\, 
        \addr_matrix_f0_0[21]\, \addr_matrix_f0_1_m_i[21]\, 
        \prdata_39_0_iv_4[22]\, \addr_matrix_f0_1_m_i[22]\, 
        \addr_matrix_f0_0_m_i[22]\, \prdata_39_0_iv_1[22]\, 
        \prdata_39_0_iv_3[22]\, \addr_data_f2_m_i[22]\, 
        \prdata_39_0_iv_2[22]\, \addr_data_f1_m_i[22]\, 
        \addr_matrix_f1[22]\, \addr_matrix_f2_m_i[22]\, 
        \prdata_39_0_iv_5[23]\, \addr_data_f3_m_i[23]\, 
        \addr_data_f2_m_i[23]\, \prdata_39_0_iv_2[23]\, 
        prdata_9_sqmuxa, \addr_data_f1_m_i[23]\, 
        \prdata_39_0_iv_1[23]\, \addr_matrix_f1[23]\, 
        \addr_matrix_f2_m_i[23]\, \prdata_39_0_iv_0[23]\, 
        \addr_matrix_f0_0[23]\, \addr_matrix_f0_1_m_i[23]\, 
        \prdata_39_0_iv_4[24]\, \addr_matrix_f0_1_m_i[24]\, 
        \addr_matrix_f0_0_m_i[24]\, \prdata_39_0_iv_1[24]\, 
        \prdata_39_0_iv_3[24]\, \addr_data_f2_m_i[24]\, 
        \prdata_39_0_iv_2[24]\, \addr_data_f1_m_i[24]\, 
        \addr_matrix_f1[24]\, \addr_matrix_f2_m_i[24]\, 
        \prdata_39_0_iv_4[25]\, \addr_matrix_f0_1_m_i[25]\, 
        \addr_matrix_f0_0_m_i[25]\, \prdata_39_0_iv_1[25]\, 
        \prdata_39_0_iv_3[25]\, \addr_data_f2_m_i[25]\, 
        \prdata_39_0_iv_2[25]\, \addr_data_f1_m_i[25]\, 
        \addr_matrix_f1[25]\, \addr_matrix_f2_m_i[25]\, 
        \prdata_39_0_iv_4[26]\, \addr_matrix_f0_1_m_i[26]\, 
        \addr_matrix_f0_0_m_i[26]\, \prdata_39_0_iv_1[26]\, 
        \prdata_39_0_iv_3[26]\, \addr_data_f2_m_i[26]\, 
        \prdata_39_0_iv_2[26]\, \addr_data_f1_m_i[26]\, 
        \addr_matrix_f1[26]\, \addr_matrix_f2_m_i[26]\, 
        \prdata_39_0_iv_4[27]\, \addr_matrix_f0_1_m_i[27]\, 
        \addr_matrix_f0_0_m_i[27]\, \prdata_39_0_iv_1[27]\, 
        \prdata_39_0_iv_3[27]\, prdata_12_sqmuxa, 
        \addr_data_f2_m_i[27]\, \prdata_39_0_iv_2[27]\, 
        \addr_data_f1_m_i[27]\, \addr_matrix_f1[27]\, 
        \addr_matrix_f2_m_i[27]\, \prdata_39_0_iv_4[28]\, 
        \addr_matrix_f0_1_m_i[28]\, \addr_matrix_f0_0_m_i[28]\, 
        \prdata_39_0_iv_1[28]\, \prdata_39_0_iv_3[28]\, 
        \addr_data_f2_m_i[28]\, \prdata_39_0_iv_2[28]\, 
        \addr_data_f1_m_i[28]\, \addr_matrix_f1[28]\, 
        \addr_matrix_f2_m_i[28]\, \prdata_39_0_iv_4[29]\, 
        \addr_matrix_f0_1_m_i[29]\, \addr_matrix_f0_0_m_i[29]\, 
        \prdata_39_0_iv_1[29]\, \prdata_39_0_iv_3[29]\, 
        \addr_data_f2_m_i[29]\, \prdata_39_0_iv_2[29]\, 
        \addr_data_f1_m_i[29]\, \addr_matrix_f1[29]\, 
        \addr_matrix_f2_m_i[29]\, \prdata_39_0_iv_4[30]\, 
        \addr_matrix_f0_1_m_i[30]\, \addr_matrix_f0_0_m_i[30]\, 
        \prdata_39_0_iv_1[30]\, \prdata_39_0_iv_3[30]\, 
        \addr_data_f2_m_i[30]\, \prdata_39_0_iv_2[30]\, 
        \addr_data_f1_m_i[30]\, \addr_matrix_f1[30]\, 
        \addr_matrix_f2_m_i[30]\, \prdata_39_0_iv_4[31]\, 
        \addr_matrix_f0_1_m_i[31]\, \addr_matrix_f0_0_m_i[31]\, 
        \prdata_39_0_iv_1[31]\, \prdata_39_0_iv_3[31]\, 
        \addr_data_f2_m_i[31]\, \prdata_39_0_iv_2[31]\, 
        \addr_data_f1_m_i[31]\, \addr_matrix_f1[31]\, 
        \addr_matrix_f2_m_i[31]\, \pirq_2_i_a2_8[15]\, 
        \pirq_2_i_a2_5[15]\, \pirq_2_i_a2_7[15]\, 
        \pirq_2_i_a2_3[15]\, \pirq_2_i_a2_6[15]\, 
        \pirq_2_i_a2_1[15]\, N_153, \status_new_err_0[3]\, N_151, 
        N_149, N_147, N_145, N_143, N_141, N_139, N_137, 
        \status_full_0[2]\, N_136, \status_full_0[1]\, N_135, 
        \status_full_0[0]\, \prdata_39[31]\, \prdata_39[30]\, 
        \prdata_39[29]\, \prdata_39[28]\, \prdata_39[27]\, 
        \prdata_39[26]\, \prdata_39[25]\, \prdata_39[24]\, 
        \prdata_39[23]\, \prdata_39[22]\, \prdata_39[21]\, 
        \prdata_39[20]\, \prdata_39[19]\, \prdata_39[18]\, 
        \prdata_39[17]\, \prdata_39[16]\, \prdata_39[15]\, 
        \prdata_39[14]\, \delta_snapshot_m_i[14]\, 
        \prdata_39[13]\, \delta_snapshot_m_i[13]\, 
        \prdata_39[11]\, \prdata_39[10]\, 
        \nb_burst_available_m_i[10]\, \prdata_39[9]\, 
        \prdata_39[8]\, \prdata_39[7]\, \prdata_39[6]\, 
        \prdata_39[5]\, \prdata_39[4]\, \prdata_39[3]\, 
        data_shaping_R0_m_i, \prdata_39[2]\, \prdata_39[1]\, 
        \prdata_39[0]\, \prdata_39[12]\, \delta_snapshot_m_i[12]\, 
        N_155_i_0, N_138, \status_full_0[3]\, 
        status_ready_matrix_f0_1, N_169, \addr_matrix_f0_0[1]\, 
        \addr_matrix_f0_1[1]\, \addr_matrix_f1[1]\, 
        \addr_matrix_f2[1]\, N_163, prdata_8_sqmuxa, 
        status_ready_matrix_f1, \addr_matrix_f0_0[2]\, 
        \addr_matrix_f0_1[2]\, \addr_matrix_f2[2]\, 
        status_ready_matrix_f2, \addr_matrix_f0_0[3]\, 
        \addr_matrix_f0_1[3]\, \addr_matrix_f2[3]\, 
        \data_shaping_R0_0\, status_error_anticipating_empty_fifo, 
        \addr_matrix_f0_0[4]\, \addr_matrix_f0_1[4]\, 
        \addr_matrix_f2[4]\, \data_shaping_R1_0\, 
        status_error_bad_component_error, \addr_matrix_f0_0[5]\, 
        \addr_matrix_f0_1[5]\, \addr_matrix_f2[5]\, 
        \addr_matrix_f0_0[6]\, \addr_matrix_f0_1[6]\, 
        \addr_matrix_f1[6]\, \addr_matrix_f2[6]\, 
        \addr_matrix_f0_0[7]\, \addr_matrix_f0_1[7]\, 
        \addr_matrix_f2[7]\, \addr_matrix_f0_1[8]\, 
        \addr_matrix_f1[8]\, \addr_matrix_f2[8]\, 
        \addr_matrix_f0_0[9]\, \addr_matrix_f0_1[9]\, 
        \addr_matrix_f2[9]\, \addr_matrix_f0_1[10]\, 
        \addr_matrix_f2[10]\, prdata_2_sqmuxa, 
        \addr_matrix_f0_0[11]\, \addr_matrix_f0_1[11]\, 
        \addr_matrix_f2[11]\, \addr_matrix_f0_1[12]\, 
        \addr_matrix_f2[12]\, \addr_matrix_f0_1[13]\, 
        \addr_matrix_f2[13]\, \addr_matrix_f0_1[14]\, 
        \addr_matrix_f2[14]\, \addr_matrix_f0_0[15]\, 
        \addr_matrix_f0_1[15]\, \addr_matrix_f2[15]\, 
        \addr_matrix_f0_0[16]\, \addr_matrix_f0_1[16]\, 
        \addr_matrix_f2[16]\, \addr_matrix_f0_0[17]\, 
        prdata_3_sqmuxa, \addr_matrix_f0_1[17]\, prdata_5_sqmuxa, 
        \addr_matrix_f2[17]\, N_161, \addr_matrix_f0_1[18]\, 
        \addr_matrix_f2[18]\, prdata_10_sqmuxa, 
        \addr_matrix_f0_0[19]\, \addr_matrix_f0_1[19]\, 
        \addr_matrix_f2[19]\, \addr_matrix_f0_0[20]\, 
        \addr_matrix_f0_1[20]\, \addr_matrix_f2[20]\, 
        \addr_matrix_f0_1[21]\, \addr_matrix_f2[21]\, 
        \addr_matrix_f0_0[22]\, \addr_matrix_f0_1[22]\, 
        \addr_matrix_f2[22]\, \addr_matrix_f0_1[23]\, 
        \addr_matrix_f2[23]\, \addr_matrix_f0_0[24]\, 
        \addr_matrix_f0_1[24]\, \addr_matrix_f2[24]\, 
        \addr_matrix_f0_0[25]\, \addr_matrix_f0_1[25]\, 
        \addr_matrix_f2[25]\, \addr_matrix_f0_0[26]\, 
        \addr_matrix_f0_1[26]\, \addr_matrix_f2[26]\, 
        \addr_matrix_f0_0[27]\, \addr_matrix_f0_1[27]\, 
        \addr_matrix_f2[27]\, \addr_matrix_f0_0[28]\, 
        \addr_matrix_f0_1[28]\, \addr_matrix_f2[28]\, 
        \addr_matrix_f0_0[29]\, \addr_matrix_f0_1[29]\, 
        \addr_matrix_f2[29]\, \addr_matrix_f0_0[30]\, 
        \addr_matrix_f0_1[30]\, \addr_matrix_f2[30]\, 
        \addr_matrix_f0_0[31]\, \addr_matrix_f0_1[31]\, 
        \addr_matrix_f2[31]\, addr_matrix_f0_0_1_sqmuxa, 
        addr_matrix_f0_1_1_sqmuxa, addr_matrix_f1_1_sqmuxa, 
        addr_matrix_f2_1_sqmuxa, addr_data_f0_1_sqmuxa, 
        addr_data_f1_1_sqmuxa, addr_data_f2_1_sqmuxa, 
        addr_data_f3_1_sqmuxa, burst_f0_1_sqmuxa, 
        delta_f2_f0_1_sqmuxa, N_164, delta_f2_f1_1_sqmuxa, 
        delta_snapshot_1_sqmuxa, nb_burst_available_1_sqmuxa, 
        N_158, nb_snapshot_param_1_sqmuxa, \status_full_ack_8[2]\, 
        \status_full_ack_8[1]\, \status_full_ack_8[0]\, 
        \status_full_5_i_o2[0]\, \status_full_RNO[0]\, 
        \status_full_RNO[1]\, \status_full_RNO[2]\, 
        \status_full_err_RNO[0]\, \status_full_err_RNO[1]\, 
        \status_full_err_RNO[2]\, \status_full_err_RNO[3]\, 
        \status_new_err_RNO[0]\, \status_new_err_RNO[1]\, 
        \status_new_err_RNO[2]\, \status_new_err_RNO[3]\, 
        status_error_anticipating_empty_fifo_1_sqmuxa, 
        config_active_interruption_onError_0_sqmuxa, 
        \addr_matrix_f2[0]\, \addr_matrix_f0_1[0]\, 
        \addr_matrix_f0_0[0]\, status_ready_matrix_f0_0, 
        \status_full_ack_8[3]\, \status_full_RNO[3]\, \enable_f3\, 
        \enable_f2\, \enable_f1\, \enable_f0\, \data_shaping_SP1\, 
        \data_shaping_SP0\, \data_shaping_BW_c\, \burst_f2\, 
        \burst_f1\, \burst_f0\, \addr_data_f1[0]\, 
        \addr_data_f1[1]\, \addr_data_f1[2]\, \addr_data_f1[3]\, 
        \addr_data_f1[4]\, \addr_data_f1[5]\, \addr_data_f1[6]\, 
        \addr_data_f1[7]\, \addr_data_f1[8]\, \addr_data_f1[9]\, 
        \addr_data_f1[10]\, \addr_data_f1[11]\, 
        \addr_data_f1[12]\, \addr_data_f1[13]\, 
        \addr_data_f1[14]\, \addr_data_f1[15]\, 
        \addr_data_f1[16]\, \addr_data_f1[17]\, 
        \addr_data_f1[18]\, \addr_data_f1[19]\, 
        \addr_data_f1[20]\, \addr_data_f1[21]\, 
        \addr_data_f1[22]\, \addr_data_f1[23]\, 
        \addr_data_f1[24]\, \addr_data_f1[25]\, 
        \addr_data_f1[26]\, \addr_data_f1[27]\, 
        \addr_data_f1[28]\, \addr_data_f1[29]\, 
        \addr_data_f1[30]\, \addr_data_f1[31]\, \addr_data_f0[0]\, 
        \addr_data_f0[1]\, \addr_data_f0[2]\, \addr_data_f0[3]\, 
        \addr_data_f0[4]\, \addr_data_f0[5]\, \addr_data_f0[6]\, 
        \addr_data_f0[7]\, \addr_data_f0[8]\, \addr_data_f0[9]\, 
        \addr_data_f0[10]\, \addr_data_f0[11]\, 
        \addr_data_f0[12]\, \addr_data_f0[13]\, 
        \addr_data_f0[14]\, \addr_data_f0[15]\, 
        \addr_data_f0[16]\, \addr_data_f0[17]\, 
        \addr_data_f0[18]\, \addr_data_f0[19]\, 
        \addr_data_f0[20]\, \addr_data_f0[21]\, 
        \addr_data_f0[22]\, \addr_data_f0[23]\, 
        \addr_data_f0[24]\, \addr_data_f0[25]\, 
        \addr_data_f0[26]\, \addr_data_f0[27]\, 
        \addr_data_f0[28]\, \addr_data_f0[29]\, 
        \addr_data_f0[30]\, \addr_data_f0[31]\, 
        \delta_snapshot[0]\, \delta_snapshot[1]\, 
        \delta_snapshot[2]\, \delta_snapshot[3]\, 
        \delta_snapshot[4]\, \delta_snapshot[5]\, 
        \delta_snapshot[6]\, \delta_snapshot[7]\, 
        \delta_snapshot[8]\, \delta_snapshot[9]\, 
        \delta_snapshot[10]\, \delta_snapshot[11]\, 
        \delta_snapshot[12]\, \delta_snapshot[13]\, 
        \delta_snapshot[14]\, \delta_snapshot[15]\, 
        \nb_snapshot_param[0]\, \nb_snapshot_param[1]\, 
        \nb_snapshot_param[2]\, \nb_snapshot_param[3]\, 
        \nb_snapshot_param[4]\, \nb_snapshot_param[5]\, 
        \nb_snapshot_param[6]\, \nb_snapshot_param[7]\, 
        \nb_snapshot_param[8]\, \nb_snapshot_param[9]\, 
        \nb_snapshot_param[10]\, \nb_burst_available[0]\, 
        \nb_burst_available[1]\, \nb_burst_available[2]\, 
        \nb_burst_available[3]\, \nb_burst_available[4]\, 
        \nb_burst_available[5]\, \nb_burst_available[6]\, 
        \nb_burst_available[7]\, \nb_burst_available[8]\, 
        \nb_burst_available[9]\, \nb_burst_available[10]\, 
        \delta_f2_f1[0]\, \delta_f2_f1[1]\, \delta_f2_f1[2]\, 
        \delta_f2_f1[3]\, \delta_f2_f1[4]\, \delta_f2_f1[5]\, 
        \delta_f2_f1[6]\, \delta_f2_f1[7]\, \delta_f2_f1[8]\, 
        \delta_f2_f1[9]\, \delta_f2_f0[0]\, \delta_f2_f0[1]\, 
        \delta_f2_f0[2]\, \delta_f2_f0[3]\, \delta_f2_f0[4]\, 
        \delta_f2_f0[5]\, \delta_f2_f0[6]\, \delta_f2_f0[7]\, 
        \delta_f2_f0[8]\, \delta_f2_f0[9]\, \addr_data_f3[0]\, 
        \addr_data_f3[1]\, \addr_data_f3[2]\, \addr_data_f3[3]\, 
        \addr_data_f3[4]\, \addr_data_f3[5]\, \addr_data_f3[6]\, 
        \addr_data_f3[7]\, \addr_data_f3[8]\, \addr_data_f3[9]\, 
        \addr_data_f3[10]\, \addr_data_f3[11]\, 
        \addr_data_f3[12]\, \addr_data_f3[13]\, 
        \addr_data_f3[14]\, \addr_data_f3[15]\, 
        \addr_data_f3[16]\, \addr_data_f3[17]\, 
        \addr_data_f3[18]\, \addr_data_f3[19]\, 
        \addr_data_f3[20]\, \addr_data_f3[21]\, 
        \addr_data_f3[22]\, \addr_data_f3[23]\, 
        \addr_data_f3[24]\, \addr_data_f3[25]\, 
        \addr_data_f3[26]\, \addr_data_f3[27]\, 
        \addr_data_f3[28]\, \addr_data_f3[29]\, 
        \addr_data_f3[30]\, \addr_data_f3[31]\, \addr_data_f2[0]\, 
        \addr_data_f2[1]\, \addr_data_f2[2]\, \addr_data_f2[3]\, 
        \addr_data_f2[4]\, \addr_data_f2[5]\, \addr_data_f2[6]\, 
        \addr_data_f2[7]\, \addr_data_f2[8]\, \addr_data_f2[9]\, 
        \addr_data_f2[10]\, \addr_data_f2[11]\, 
        \addr_data_f2[12]\, \addr_data_f2[13]\, 
        \addr_data_f2[14]\, \addr_data_f2[15]\, 
        \addr_data_f2[16]\, \addr_data_f2[17]\, 
        \addr_data_f2[18]\, \addr_data_f2[19]\, 
        \addr_data_f2[20]\, \addr_data_f2[21]\, 
        \addr_data_f2[22]\, \addr_data_f2[23]\, 
        \addr_data_f2[24]\, \addr_data_f2[25]\, 
        \addr_data_f2[26]\, \addr_data_f2[27]\, 
        \addr_data_f2[28]\, \addr_data_f2[29]\, 
        \addr_data_f2[30]\, \addr_data_f2[31]\, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 

    addr_data_f2(31) <= \addr_data_f2[31]\;
    addr_data_f2(30) <= \addr_data_f2[30]\;
    addr_data_f2(29) <= \addr_data_f2[29]\;
    addr_data_f2(28) <= \addr_data_f2[28]\;
    addr_data_f2(27) <= \addr_data_f2[27]\;
    addr_data_f2(26) <= \addr_data_f2[26]\;
    addr_data_f2(25) <= \addr_data_f2[25]\;
    addr_data_f2(24) <= \addr_data_f2[24]\;
    addr_data_f2(23) <= \addr_data_f2[23]\;
    addr_data_f2(22) <= \addr_data_f2[22]\;
    addr_data_f2(21) <= \addr_data_f2[21]\;
    addr_data_f2(20) <= \addr_data_f2[20]\;
    addr_data_f2(19) <= \addr_data_f2[19]\;
    addr_data_f2(18) <= \addr_data_f2[18]\;
    addr_data_f2(17) <= \addr_data_f2[17]\;
    addr_data_f2(16) <= \addr_data_f2[16]\;
    addr_data_f2(15) <= \addr_data_f2[15]\;
    addr_data_f2(14) <= \addr_data_f2[14]\;
    addr_data_f2(13) <= \addr_data_f2[13]\;
    addr_data_f2(12) <= \addr_data_f2[12]\;
    addr_data_f2(11) <= \addr_data_f2[11]\;
    addr_data_f2(10) <= \addr_data_f2[10]\;
    addr_data_f2(9) <= \addr_data_f2[9]\;
    addr_data_f2(8) <= \addr_data_f2[8]\;
    addr_data_f2(7) <= \addr_data_f2[7]\;
    addr_data_f2(6) <= \addr_data_f2[6]\;
    addr_data_f2(5) <= \addr_data_f2[5]\;
    addr_data_f2(4) <= \addr_data_f2[4]\;
    addr_data_f2(3) <= \addr_data_f2[3]\;
    addr_data_f2(2) <= \addr_data_f2[2]\;
    addr_data_f2(1) <= \addr_data_f2[1]\;
    addr_data_f2(0) <= \addr_data_f2[0]\;
    addr_data_f3(31) <= \addr_data_f3[31]\;
    addr_data_f3(30) <= \addr_data_f3[30]\;
    addr_data_f3(29) <= \addr_data_f3[29]\;
    addr_data_f3(28) <= \addr_data_f3[28]\;
    addr_data_f3(27) <= \addr_data_f3[27]\;
    addr_data_f3(26) <= \addr_data_f3[26]\;
    addr_data_f3(25) <= \addr_data_f3[25]\;
    addr_data_f3(24) <= \addr_data_f3[24]\;
    addr_data_f3(23) <= \addr_data_f3[23]\;
    addr_data_f3(22) <= \addr_data_f3[22]\;
    addr_data_f3(21) <= \addr_data_f3[21]\;
    addr_data_f3(20) <= \addr_data_f3[20]\;
    addr_data_f3(19) <= \addr_data_f3[19]\;
    addr_data_f3(18) <= \addr_data_f3[18]\;
    addr_data_f3(17) <= \addr_data_f3[17]\;
    addr_data_f3(16) <= \addr_data_f3[16]\;
    addr_data_f3(15) <= \addr_data_f3[15]\;
    addr_data_f3(14) <= \addr_data_f3[14]\;
    addr_data_f3(13) <= \addr_data_f3[13]\;
    addr_data_f3(12) <= \addr_data_f3[12]\;
    addr_data_f3(11) <= \addr_data_f3[11]\;
    addr_data_f3(10) <= \addr_data_f3[10]\;
    addr_data_f3(9) <= \addr_data_f3[9]\;
    addr_data_f3(8) <= \addr_data_f3[8]\;
    addr_data_f3(7) <= \addr_data_f3[7]\;
    addr_data_f3(6) <= \addr_data_f3[6]\;
    addr_data_f3(5) <= \addr_data_f3[5]\;
    addr_data_f3(4) <= \addr_data_f3[4]\;
    addr_data_f3(3) <= \addr_data_f3[3]\;
    addr_data_f3(2) <= \addr_data_f3[2]\;
    addr_data_f3(1) <= \addr_data_f3[1]\;
    addr_data_f3(0) <= \addr_data_f3[0]\;
    nb_burst_available(10) <= \nb_burst_available[10]\;
    nb_burst_available(9) <= \nb_burst_available[9]\;
    nb_burst_available(8) <= \nb_burst_available[8]\;
    nb_burst_available(7) <= \nb_burst_available[7]\;
    nb_burst_available(6) <= \nb_burst_available[6]\;
    nb_burst_available(5) <= \nb_burst_available[5]\;
    nb_burst_available(4) <= \nb_burst_available[4]\;
    nb_burst_available(3) <= \nb_burst_available[3]\;
    nb_burst_available(2) <= \nb_burst_available[2]\;
    nb_burst_available(1) <= \nb_burst_available[1]\;
    nb_burst_available(0) <= \nb_burst_available[0]\;
    addr_data_f1(31) <= \addr_data_f1[31]\;
    addr_data_f1(30) <= \addr_data_f1[30]\;
    addr_data_f1(29) <= \addr_data_f1[29]\;
    addr_data_f1(28) <= \addr_data_f1[28]\;
    addr_data_f1(27) <= \addr_data_f1[27]\;
    addr_data_f1(26) <= \addr_data_f1[26]\;
    addr_data_f1(25) <= \addr_data_f1[25]\;
    addr_data_f1(24) <= \addr_data_f1[24]\;
    addr_data_f1(23) <= \addr_data_f1[23]\;
    addr_data_f1(22) <= \addr_data_f1[22]\;
    addr_data_f1(21) <= \addr_data_f1[21]\;
    addr_data_f1(20) <= \addr_data_f1[20]\;
    addr_data_f1(19) <= \addr_data_f1[19]\;
    addr_data_f1(18) <= \addr_data_f1[18]\;
    addr_data_f1(17) <= \addr_data_f1[17]\;
    addr_data_f1(16) <= \addr_data_f1[16]\;
    addr_data_f1(15) <= \addr_data_f1[15]\;
    addr_data_f1(14) <= \addr_data_f1[14]\;
    addr_data_f1(13) <= \addr_data_f1[13]\;
    addr_data_f1(12) <= \addr_data_f1[12]\;
    addr_data_f1(11) <= \addr_data_f1[11]\;
    addr_data_f1(10) <= \addr_data_f1[10]\;
    addr_data_f1(9) <= \addr_data_f1[9]\;
    addr_data_f1(8) <= \addr_data_f1[8]\;
    addr_data_f1(7) <= \addr_data_f1[7]\;
    addr_data_f1(6) <= \addr_data_f1[6]\;
    addr_data_f1(5) <= \addr_data_f1[5]\;
    addr_data_f1(4) <= \addr_data_f1[4]\;
    addr_data_f1(3) <= \addr_data_f1[3]\;
    addr_data_f1(2) <= \addr_data_f1[2]\;
    addr_data_f1(1) <= \addr_data_f1[1]\;
    addr_data_f1(0) <= \addr_data_f1[0]\;
    delta_f2_f1(9) <= \delta_f2_f1[9]\;
    delta_f2_f1(8) <= \delta_f2_f1[8]\;
    delta_f2_f1(7) <= \delta_f2_f1[7]\;
    delta_f2_f1(6) <= \delta_f2_f1[6]\;
    delta_f2_f1(5) <= \delta_f2_f1[5]\;
    delta_f2_f1(4) <= \delta_f2_f1[4]\;
    delta_f2_f1(3) <= \delta_f2_f1[3]\;
    delta_f2_f1(2) <= \delta_f2_f1[2]\;
    delta_f2_f1(1) <= \delta_f2_f1[1]\;
    delta_f2_f1(0) <= \delta_f2_f1[0]\;
    addr_data_f0(31) <= \addr_data_f0[31]\;
    addr_data_f0(30) <= \addr_data_f0[30]\;
    addr_data_f0(29) <= \addr_data_f0[29]\;
    addr_data_f0(28) <= \addr_data_f0[28]\;
    addr_data_f0(27) <= \addr_data_f0[27]\;
    addr_data_f0(26) <= \addr_data_f0[26]\;
    addr_data_f0(25) <= \addr_data_f0[25]\;
    addr_data_f0(24) <= \addr_data_f0[24]\;
    addr_data_f0(23) <= \addr_data_f0[23]\;
    addr_data_f0(22) <= \addr_data_f0[22]\;
    addr_data_f0(21) <= \addr_data_f0[21]\;
    addr_data_f0(20) <= \addr_data_f0[20]\;
    addr_data_f0(19) <= \addr_data_f0[19]\;
    addr_data_f0(18) <= \addr_data_f0[18]\;
    addr_data_f0(17) <= \addr_data_f0[17]\;
    addr_data_f0(16) <= \addr_data_f0[16]\;
    addr_data_f0(15) <= \addr_data_f0[15]\;
    addr_data_f0(14) <= \addr_data_f0[14]\;
    addr_data_f0(13) <= \addr_data_f0[13]\;
    addr_data_f0(12) <= \addr_data_f0[12]\;
    addr_data_f0(11) <= \addr_data_f0[11]\;
    addr_data_f0(10) <= \addr_data_f0[10]\;
    addr_data_f0(9) <= \addr_data_f0[9]\;
    addr_data_f0(8) <= \addr_data_f0[8]\;
    addr_data_f0(7) <= \addr_data_f0[7]\;
    addr_data_f0(6) <= \addr_data_f0[6]\;
    addr_data_f0(5) <= \addr_data_f0[5]\;
    addr_data_f0(4) <= \addr_data_f0[4]\;
    addr_data_f0(3) <= \addr_data_f0[3]\;
    addr_data_f0(2) <= \addr_data_f0[2]\;
    addr_data_f0(1) <= \addr_data_f0[1]\;
    addr_data_f0(0) <= \addr_data_f0[0]\;
    delta_f2_f0(9) <= \delta_f2_f0[9]\;
    delta_f2_f0(8) <= \delta_f2_f0[8]\;
    delta_f2_f0(7) <= \delta_f2_f0[7]\;
    delta_f2_f0(6) <= \delta_f2_f0[6]\;
    delta_f2_f0(5) <= \delta_f2_f0[5]\;
    delta_f2_f0(4) <= \delta_f2_f0[4]\;
    delta_f2_f0(3) <= \delta_f2_f0[3]\;
    delta_f2_f0(2) <= \delta_f2_f0[2]\;
    delta_f2_f0(1) <= \delta_f2_f0[1]\;
    delta_f2_f0(0) <= \delta_f2_f0[0]\;
    delta_snapshot(15) <= \delta_snapshot[15]\;
    delta_snapshot(14) <= \delta_snapshot[14]\;
    delta_snapshot(13) <= \delta_snapshot[13]\;
    delta_snapshot(12) <= \delta_snapshot[12]\;
    delta_snapshot(11) <= \delta_snapshot[11]\;
    delta_snapshot(10) <= \delta_snapshot[10]\;
    delta_snapshot(9) <= \delta_snapshot[9]\;
    delta_snapshot(8) <= \delta_snapshot[8]\;
    delta_snapshot(7) <= \delta_snapshot[7]\;
    delta_snapshot(6) <= \delta_snapshot[6]\;
    delta_snapshot(5) <= \delta_snapshot[5]\;
    delta_snapshot(4) <= \delta_snapshot[4]\;
    delta_snapshot(3) <= \delta_snapshot[3]\;
    delta_snapshot(2) <= \delta_snapshot[2]\;
    delta_snapshot(1) <= \delta_snapshot[1]\;
    delta_snapshot(0) <= \delta_snapshot[0]\;
    nb_snapshot_param(10) <= \nb_snapshot_param[10]\;
    nb_snapshot_param(9) <= \nb_snapshot_param[9]\;
    nb_snapshot_param(8) <= \nb_snapshot_param[8]\;
    nb_snapshot_param(7) <= \nb_snapshot_param[7]\;
    nb_snapshot_param(6) <= \nb_snapshot_param[6]\;
    nb_snapshot_param(5) <= \nb_snapshot_param[5]\;
    nb_snapshot_param(4) <= \nb_snapshot_param[4]\;
    nb_snapshot_param(3) <= \nb_snapshot_param[3]\;
    nb_snapshot_param(2) <= \nb_snapshot_param[2]\;
    nb_snapshot_param(1) <= \nb_snapshot_param[1]\;
    nb_snapshot_param(0) <= \nb_snapshot_param[0]\;
    enable_f0 <= \enable_f0\;
    data_shaping_BW_c <= \data_shaping_BW_c\;
    burst_f2 <= \burst_f2\;
    burst_f1 <= \burst_f1\;
    burst_f0 <= \burst_f0\;
    enable_f3 <= \enable_f3\;
    enable_f2 <= \enable_f2\;
    data_shaping_SP1 <= \data_shaping_SP1\;
    enable_f1 <= \enable_f1\;
    data_shaping_SP0 <= \data_shaping_SP0\;
    data_shaping_R1_0 <= \data_shaping_R1_0\;
    data_shaping_R0_0 <= \data_shaping_R0_0\;

    \prdata_RNO_7[29]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[29]\, C
         => \addr_matrix_f2_m_i[29]\, Y => \prdata_39_0_iv_1[29]\);
    
    \reg_wp.addr_data_f3[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[17]\);
    
    \reg_wp.delta_f2_f1[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[1]\);
    
    \reg_sp.addr_matrix_f1[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[6]\);
    
    \prdata_RNO_5[14]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[14]\, C => \addr_matrix_f0_1_m_i[14]\, 
        Y => \prdata_39_0_iv_0[14]\);
    
    \prdata_RNO_2[14]\ : NOR3C
      port map(A => \prdata_39_0_iv_1[14]\, B => 
        \prdata_39_0_iv_0[14]\, C => \prdata_39_0_iv_3[14]\, Y
         => \prdata_39_0_iv_6[14]\);
    
    \reg_sp.addr_matrix_f0_0[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[2]\);
    
    \reg_wp.addr_data_f3[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[25]\);
    
    \prdata_RNO_0[8]\ : NOR3C
      port map(A => \prdata_39_0_iv_0[8]\, B => 
        \delta_f2_f1_m_i[8]\, C => \prdata_39_0_iv_6[8]\, Y => 
        \prdata_39_0_iv_9[8]\);
    
    \reg_wp.addr_data_f3[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[26]\);
    
    \reg_wp.nb_snapshot_param[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[2]\);
    
    \reg_wp.delta_f2_f0[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[2]\);
    
    \reg_wp.addr_data_f3_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_168, B => N_157, C => un1_apbi_2, Y => 
        addr_data_f3_1_sqmuxa);
    
    \prdata_RNO_5[7]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[7]\, B => 
        \addr_matrix_f0_0_m_i[7]\, C => \delta_f2_f1_m_i[7]\, Y
         => \prdata_39_0_iv_5[7]\);
    
    \reg_wp.addr_data_f2[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[29]\);
    
    prdata_18_sqmuxa_0_a2 : NOR3C
      port map(A => N_158, B => N_159, C => apbi_c_19, Y => 
        prdata_18_sqmuxa);
    
    \reg_sp.addr_matrix_f0_1[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[22]\);
    
    \prdata_RNO_7[3]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[3]\, B => 
        \addr_matrix_f0_0_m_i[3]\, C => \status_full_m_i[3]\, Y
         => \prdata_39_0_iv_6[3]\);
    
    \prdata_RNO_8[28]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[28]\, Y
         => \addr_matrix_f2_m_i[28]\);
    
    \prdata_RNO_6[1]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[1]\, C
         => enable_f1_m_i, Y => \prdata_39_0_iv_8[1]\);
    
    \prdata_RNO_4[29]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[29]\, Y
         => \addr_data_f1_m_i[29]\);
    
    \reg_wp.nb_snapshot_param[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[9]\);
    
    \reg_wp.nb_burst_available[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[7]\);
    
    \prdata_RNO[8]\ : OR3C
      port map(A => \prdata_39_0_iv_9[8]\, B => 
        \prdata_39_0_iv_8[8]\, C => \prdata_39_0_iv_10[8]\, Y => 
        \prdata_39[8]\);
    
    \prdata_RNO_1[13]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[13]\, 
        Y => \delta_snapshot_m_i[13]\);
    
    \prdata_RNO_6[18]\ : OR3C
      port map(A => N_161, B => N_168_0, C => \addr_data_f2[18]\, 
        Y => \addr_data_f2_m_i[18]\);
    
    \prdata[26]\ : DFN1C0
      port map(D => \prdata_39[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(26));
    
    \prdata_RNO_19[0]\ : AOI1B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[0]\, C
         => data_shaping_BW_m_i, Y => \prdata_39_0_iv_5[0]\);
    
    \reg_sp.addr_matrix_f0_0[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[4]\);
    
    \prdata_RNO_0[29]\ : AOI1B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[29]\, C
         => \addr_data_f2_m_i[29]\, Y => \prdata_39_0_iv_3[29]\);
    
    \reg_wp.delta_f2_f0_1_sqmuxa_0_a2_2\ : NOR3B
      port map(A => apbi_c_0, B => apbi_c_23, C => apbi_c_24, Y
         => N_158);
    
    \reg_wp.addr_data_f0_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_930, B => apbi_c_21, C => N_931, Y => 
        addr_data_f0_1_sqmuxa);
    
    \prdata_RNO_7[10]\ : OR2B
      port map(A => \nb_snapshot_param[10]\, B => 
        prdata_18_sqmuxa, Y => \nb_snapshot_param_m_i[10]\);
    
    \reg_wp.addr_data_f2[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[13]\);
    
    \reg_wp.addr_data_f2[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[10]\);
    
    \reg_sp.addr_matrix_f0_1[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[2]\);
    
    \reg_wp.addr_data_f3[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[2]\);
    
    \reg_wp.addr_data_f3_1_sqmuxa_0_a2_0\ : NOR3A
      port map(A => N_168, B => N_157, C => un1_apbi_2, Y => 
        addr_data_f3_1_sqmuxa_0);
    
    \reg_sp.addr_matrix_f0_1[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[1]\);
    
    \prdata_RNO_11[1]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[1]\, Y
         => \addr_data_f1_m_i[1]\);
    
    \apbo.pirq_RNO_4[15]\ : NOR2
      port map(A => status_new_err_0_2, B => status_new_err_3, Y
         => \pirq_2_i_a2_1[15]\);
    
    \prdata_RNO_4[14]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[14]\, 
        C => \addr_matrix_f2_m_i[14]\, Y => 
        \prdata_39_0_iv_1[14]\);
    
    \reg_sp.addr_matrix_f0_0[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[31]\);
    
    \prdata_RNO_13[6]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[6]\, Y
         => \delta_f2_f1_m_i[6]\);
    
    \prdata_RNO_16[6]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[6]\, Y
         => \delta_f2_f0_m_i[6]\);
    
    \reg_sp.addr_matrix_f0_1[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[19]\);
    
    \reg_sp.status_ready_matrix_f2\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_ready_matrix_f2);
    
    \prdata_RNO_6[20]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[20]\, 
        Y => \addr_matrix_f0_0_m_i[20]\);
    
    \reg_wp.addr_data_f0[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[8]\);
    
    \prdata_RNO_6[4]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[4]\, B => 
        \addr_matrix_f0_0_m_i[4]\, C => \prdata_39_0_iv_1[4]\, Y
         => \prdata_39_0_iv_6[4]\);
    
    \prdata_RNO_6[31]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[31]\, 
        Y => \addr_matrix_f0_0_m_i[31]\);
    
    \apbo.pirq_RNO_0[15]\ : NOR3A
      port map(A => \pirq_2_i_a2_3[15]\, B => 
        status_full_err_0(1), C => status_full_err_0(0), Y => 
        \pirq_2_i_a2_7[15]\);
    
    \reg_sp.addr_matrix_f0_1[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[9]\);
    
    \prdata_RNO_3[6]\ : NOR3C
      port map(A => \addr_matrix_f2_m_i[6]\, B => 
        \addr_matrix_f1_m_i[6]\, C => \delta_snapshot_m_i[6]\, Y
         => \prdata_39_0_iv_6[6]\);
    
    \prdata_RNO_18[1]\ : OR2B
      port map(A => \status_full_0[1]\, B => prdata_13_sqmuxa, Y
         => \status_full_m_i[1]\);
    
    \reg_wp.delta_snapshot_1_sqmuxa_0_o2_0\ : OR3C
      port map(A => apbi_c_22, B => N_928, C => apbi_c_20, Y => 
        N_931);
    
    \reg_sp.addr_matrix_f0_0[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[24]\);
    
    \prdata_RNO_11[10]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[10]\, Y
         => \addr_data_f0_m_i[10]\);
    
    \reg_wp.addr_data_f2[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[11]\);
    
    \reg_sp.addr_matrix_f0_0[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[25]\);
    
    \reg_sp.addr_matrix_f0_0[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[16]\);
    
    \prdata_RNO_9[6]\ : OR2B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[6]\, Y
         => \addr_matrix_f1_m_i[6]\);
    
    \reg_sp.addr_matrix_f0_1_1_sqmuxa_0_a2_0\ : NOR2A
      port map(A => apbi_c_19, B => un1_apbi_2, Y => N_166);
    
    \prdata_RNO_9[7]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[7]\, C
         => \addr_data_f2_m_i[7]\, Y => \prdata_39_0_iv_3[7]\);
    
    \prdata_RNO_8[0]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[0]\, C
         => \addr_data_f1_m_i[0]\, Y => \prdata_39_0_iv_3[0]\);
    
    \prdata_RNO_16[9]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[9]\, 
        Y => \addr_data_f2_m_i[9]\);
    
    \prdata_RNO[7]\ : OR3C
      port map(A => \prdata_39_0_iv_9[7]\, B => 
        \prdata_39_0_iv_8[7]\, C => \prdata_39_0_iv_10[7]\, Y => 
        \prdata_39[7]\);
    
    \prdata_RNO_5[13]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[13]\, C => \addr_matrix_f0_1_m_i[13]\, 
        Y => \prdata_39_0_iv_0[13]\);
    
    \prdata_RNO_2[13]\ : NOR3C
      port map(A => \prdata_39_0_iv_1[13]\, B => 
        \prdata_39_0_iv_0[13]\, C => \prdata_39_0_iv_3[13]\, Y
         => \prdata_39_0_iv_6[13]\);
    
    prdata_16_sqmuxa_0_a2 : NOR2A
      port map(A => N_164, B => N_157, Y => prdata_16_sqmuxa);
    
    \prdata_RNO_7[1]\ : NOR3C
      port map(A => \addr_matrix_f2_m_i[1]\, B => 
        \addr_matrix_f1_m_i[1]\, C => \prdata_39_0_iv_2[1]\, Y
         => \prdata_39_0_iv_7[1]\);
    
    \reg_wp.addr_data_f3[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[5]\);
    
    \prdata_RNO_9[15]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[15]\, 
        Y => \delta_snapshot_m_i[15]\);
    
    \prdata_RNO_7[25]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[25]\, C
         => \addr_matrix_f2_m_i[25]\, Y => \prdata_39_0_iv_1[25]\);
    
    \prdata_RNO_10[2]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[2]\, 
        Y => \addr_data_f2_m_i[2]\);
    
    \reg_wp.addr_data_f3[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[22]\);
    
    \reg_wp.status_new_err_RNO_0[3]\ : NOR3A
      port map(A => N_933_0, B => \status_new_err_0[3]\, C => 
        status_new_err_3, Y => N_153);
    
    \prdata_RNO_8[27]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[27]\, Y
         => \addr_matrix_f2_m_i[27]\);
    
    \reg_sp.addr_matrix_f0_1[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[4]\);
    
    \reg_wp.burst_f2\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \burst_f2\);
    
    \reg_sp.addr_matrix_f1[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[0]\);
    
    \prdata_RNO_11[7]\ : OR2B
      port map(A => \nb_burst_available[7]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[7]\);
    
    \reg_wp.status_full_err[3]\ : DFN1C0
      port map(D => \status_full_err_RNO[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_full_err[3]\);
    
    \prdata_RNO_20[1]\ : OR3A
      port map(A => status_ready_matrix_f0_1, B => N_157, C => 
        N_169, Y => status_ready_matrix_f0_1_m_i);
    
    \prdata_RNO_19[4]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[4]\, 
        Y => \addr_matrix_f2_m_i[4]\);
    
    \prdata_RNO_2[24]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[24]\, B => 
        \addr_matrix_f0_0_m_i[24]\, C => \prdata_39_0_iv_1[24]\, 
        Y => \prdata_39_0_iv_4[24]\);
    
    \prdata_RNO_8[4]\ : NOR3C
      port map(A => \addr_data_f3_m_i[4]\, B => 
        \addr_data_f2_m_i[4]\, C => \prdata_39_0_iv_5[4]\, Y => 
        \prdata_39_0_iv_9[4]\);
    
    \prdata_RNO[18]\ : OR3C
      port map(A => \prdata_39_0_iv_1[18]\, B => 
        \prdata_39_0_iv_0[18]\, C => \prdata_39_0_iv_5[18]\, Y
         => \prdata_39[18]\);
    
    \status_full_ack[1]\ : DFN1C0
      port map(D => \status_full_ack_8[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => status_full_ack(1));
    
    \prdata_RNO_1[30]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[30]\, C
         => \addr_data_f1_m_i[30]\, Y => \prdata_39_0_iv_2[30]\);
    
    \reg_sp.addr_matrix_f0_0_1_sqmuxa_0_o2\ : NOR2
      port map(A => un1_apbi_2, B => apbi_c_19, Y => N_930);
    
    \prdata_RNO_6[17]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[17]\, 
        Y => \addr_matrix_f0_0_m_i[17]\);
    
    \reg_sp.addr_matrix_f1[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[8]\);
    
    \prdata_RNO_4[25]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[25]\, Y
         => \addr_data_f1_m_i[25]\);
    
    \prdata_RNO_1[3]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[3]\, B => 
        \prdata_39_0_iv_2[3]\, C => \prdata_39_0_iv_9[3]\, Y => 
        \prdata_39_0_iv_12[3]\);
    
    \prdata_RNO_16[8]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[8]\, 
        Y => \addr_data_f2_m_i[8]\);
    
    \prdata_RNO_5[21]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[21]\, Y
         => \addr_data_f3_m_i[21]\);
    
    \prdata_RNO_5[26]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[26]\, 
        Y => \addr_matrix_f0_1_m_i[26]\);
    
    prdata_0_sqmuxa_0_a2_0 : NOR2
      port map(A => apbi_c_20, B => apbi_c_19, Y => N_161);
    
    \prdata[7]\ : DFN1C0
      port map(D => \prdata_39[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(7));
    
    \reg_sp.config_active_interruption_onError\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => config_active_interruption_onError_0_sqmuxa, Q => 
        config_active_interruption_onError);
    
    \prdata_RNO_3[19]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[19]\, Y
         => \addr_data_f2_m_i[19]\);
    
    \prdata_RNO_4[5]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \burst_f1\, Y => 
        burst_f1_m_i);
    
    \prdata_RNO_7[28]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[28]\, C
         => \addr_matrix_f2_m_i[28]\, Y => \prdata_39_0_iv_1[28]\);
    
    \reg_wp.delta_f2_f1[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[7]\);
    
    \prdata_RNO_12[0]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[0]\, 
        Y => \addr_matrix_f0_1_m_i[0]\);
    
    \prdata_RNO_0[25]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[25]\, 
        C => \addr_data_f2_m_i[25]\, Y => \prdata_39_0_iv_3[25]\);
    
    \prdata[14]\ : DFN1C0
      port map(D => \prdata_39[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(14));
    
    \prdata_RNO_11[3]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[3]\, Y
         => \delta_f2_f0_m_i[3]\);
    
    \prdata_RNO_4[13]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[13]\, 
        C => \addr_matrix_f2_m_i[13]\, Y => 
        \prdata_39_0_iv_1[13]\);
    
    \prdata_RNO_2[9]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[9]\, B => 
        \prdata_39_0_iv_2[9]\, C => \nb_burst_available_m_i[9]\, 
        Y => \prdata_39_0_iv_10[9]\);
    
    prdata_12_sqmuxa_0_a2_0 : NOR2A
      port map(A => N_168, B => N_157, Y => prdata_12_sqmuxa_0);
    
    \reg_wp.status_full_RNO_0[2]\ : NOR3A
      port map(A => N_933_0, B => \status_full_0[2]\, C => 
        status_full(2), Y => N_137);
    
    \prdata_RNO_12[4]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[4]\, 
        Y => \addr_matrix_f0_1_m_i[4]\);
    
    \prdata_RNO_5[22]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[22]\, 
        Y => \addr_matrix_f0_1_m_i[22]\);
    
    \reg_wp.addr_data_f2[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[15]\);
    
    \reg_wp.addr_data_f2[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[16]\);
    
    \reg_sp.config_active_interruption_onError_0_sqmuxa_0_a2\ : 
        NOR3A
      port map(A => N_930, B => apbi_c_20, C => N_169, Y => 
        config_active_interruption_onError_0_sqmuxa);
    
    \reg_sp.addr_matrix_f2[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[15]\);
    
    \prdata_RNO[23]\ : OR3C
      port map(A => \prdata_39_0_iv_1[23]\, B => 
        \prdata_39_0_iv_0[23]\, C => \prdata_39_0_iv_5[23]\, Y
         => \prdata_39[23]\);
    
    \reg_wp.burst_f0_1_sqmuxa_0_a2\ : NOR3
      port map(A => N_157, B => un1_apbi_2, C => N_163, Y => 
        burst_f0_1_sqmuxa);
    
    \reg_wp.addr_data_f0[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[7]\);
    
    \reg_sp.addr_matrix_f0_0[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[10]\);
    
    \prdata_RNO_6[0]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[0]\, B => 
        \addr_matrix_f0_0_m_i[0]\, C => \prdata_39_0_iv_1[0]\, Y
         => \prdata_39_0_iv_7[0]\);
    
    \reg_wp.addr_data_f1[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[27]\);
    
    \reg_wp.nb_burst_available[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[9]\);
    
    \reg_wp.addr_data_f1[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[8]\);
    
    \prdata_RNO_4[28]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[28]\, Y
         => \addr_data_f1_m_i[28]\);
    
    \reg_sp.addr_matrix_f0_0[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[13]\);
    
    \apbo.pirq_RNO[15]\ : OR3C
      port map(A => \pirq_2_i_a2_7[15]\, B => \pirq_2_i_a2_6[15]\, 
        C => \pirq_2_i_a2_8[15]\, Y => N_155_i_0);
    
    \reg_sp.addr_matrix_f2[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[12]\);
    
    \prdata_RNO_1[10]\ : OR2B
      port map(A => \nb_burst_available[10]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[10]\);
    
    \reg_sp.config_active_interruption_onError_0_sqmuxa_0_a2_0\ : 
        OR3A
      port map(A => N_928, B => apbi_c_21, C => apbi_c_22, Y => 
        N_169);
    
    \reg_wp.addr_data_f1[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[5]\);
    
    \prdata_RNO_3[21]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[21]\, Y
         => \addr_matrix_f2_m_i[21]\);
    
    \prdata_RNO_15[3]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[3]\, 
        Y => \addr_matrix_f0_0_m_i[3]\);
    
    \prdata_RNO_3[26]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[26]\, Y
         => \addr_data_f2_m_i[26]\);
    
    \prdata_RNO_8[19]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[19]\, Y
         => \addr_matrix_f2_m_i[19]\);
    
    \prdata_RNO_3[1]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[1]\, C
         => \addr_data_f2_m_i[1]\, Y => \prdata_39_0_iv_4[1]\);
    
    \prdata_RNO_20[0]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[0]\, Y
         => \addr_matrix_f2_m_i[0]\);
    
    \prdata[27]\ : DFN1C0
      port map(D => \prdata_39[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(27));
    
    \prdata_RNO[12]\ : OR3C
      port map(A => \prdata_39_0_iv_2[12]\, B => 
        \delta_snapshot_m_i[12]\, C => \prdata_39_0_iv_6[12]\, Y
         => \prdata_39[12]\);
    
    \reg_sp.addr_matrix_f2[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[17]\);
    
    \reg_wp.addr_data_f2[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[4]\);
    
    \prdata_RNO_2[3]\ : NOR3C
      port map(A => \nb_snapshot_param_m_i[3]\, B => 
        \prdata_39_0_iv_6[3]\, C => \prdata_39_0_iv_11[3]\, Y => 
        \prdata_39_0_iv_13[3]\);
    
    \prdata_RNO_15[4]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[4]\, Y
         => \addr_data_f3_m_i[4]\);
    
    \prdata[28]\ : DFN1C0
      port map(D => \prdata_39[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(28));
    
    \prdata_RNO_0[28]\ : AOI1B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[28]\, C
         => \addr_data_f2_m_i[28]\, Y => \prdata_39_0_iv_3[28]\);
    
    \reg_wp.addr_data_f3[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[13]\);
    
    \prdata_RNO_2[23]\ : NOR3C
      port map(A => \addr_data_f3_m_i[23]\, B => 
        \addr_data_f2_m_i[23]\, C => \prdata_39_0_iv_2[23]\, Y
         => \prdata_39_0_iv_5[23]\);
    
    \reg_sp.addr_matrix_f2[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[25]\);
    
    \reg_wp.addr_data_f3[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[10]\);
    
    \prdata_RNO_9[8]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[8]\, C
         => \addr_data_f2_m_i[8]\, Y => \prdata_39_0_iv_3[8]\);
    
    \prdata_RNO_13[0]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[0]\, 
        Y => \addr_matrix_f0_0_m_i[0]\);
    
    \reg_wp.data_shaping_R0\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => data_shaping_R0);
    
    \reg_wp.addr_data_f2[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[6]\);
    
    \prdata_RNO_14[7]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[7]\, 
        Y => \addr_matrix_f0_0_m_i[7]\);
    
    \prdata_RNO[24]\ : OR3C
      port map(A => \prdata_39_0_iv_3[24]\, B => 
        \prdata_39_0_iv_2[24]\, C => \prdata_39_0_iv_4[24]\, Y
         => \prdata_39[24]\);
    
    \prdata_RNO_7[0]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[0]\, C
         => \addr_data_f2_m_i[0]\, Y => \prdata_39_0_iv_4[0]\);
    
    \prdata_RNO[10]\ : OR3C
      port map(A => \prdata_39_0_iv_7[10]\, B => 
        \nb_burst_available_m_i[10]\, C => \prdata_39_0_iv_8[10]\, 
        Y => \prdata_39[10]\);
    
    \reg_sp.addr_matrix_f0_1[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[17]\);
    
    \reg_wp.data_shaping_SP1\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => \data_shaping_SP1\);
    
    \reg_sp.addr_matrix_f2[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[22]\);
    
    \prdata_RNO_3[22]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[22]\, Y
         => \addr_data_f2_m_i[22]\);
    
    \reg_wp.status_full_err_RNO[1]\ : OA1B
      port map(A => apbi_c_55, B => \status_full_5_i_o2[0]\, C
         => N_141, Y => \status_full_err_RNO[1]\);
    
    \reg_wp.delta_snapshot[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[1]\);
    
    \reg_sp.addr_matrix_f0_1[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[21]\);
    
    prdata_2_sqmuxa_0_a2_0 : NOR3B
      port map(A => N_159, B => N_928, C => apbi_c_19, Y => 
        prdata_2_sqmuxa_0);
    
    \prdata_RNO_0[11]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[11]\, 
        C => \prdata_39_0_iv_1[11]\, Y => \prdata_39_0_iv_5[11]\);
    
    \prdata_RNO_7[27]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[27]\, C
         => \addr_matrix_f2_m_i[27]\, Y => \prdata_39_0_iv_1[27]\);
    
    \prdata_RNO_0[16]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[16]\, 
        C => \addr_data_f2_m_i[16]\, Y => \prdata_39_0_iv_3[16]\);
    
    \reg_wp.addr_data_f3[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[11]\);
    
    \reg_sp.addr_matrix_f2[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[27]\);
    
    \reg_sp.addr_matrix_f1[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[29]\);
    
    \reg_wp.delta_f2_f0[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[1]\);
    
    \reg_wp.burst_f0_1_sqmuxa_0_a2_0\ : OR3B
      port map(A => apbi_c_22, B => N_928, C => apbi_c_21, Y => 
        N_163);
    
    \reg_wp.addr_data_f1[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[17]\);
    
    \reg_wp.status_new_err_RNO[3]\ : OA1B
      port map(A => apbi_c_61, B => \status_full_5_i_o2[0]\, C
         => N_153, Y => \status_new_err_RNO[3]\);
    
    \prdata_RNO_6[6]\ : AOI1B
      port map(A => \status_full_err[2]\, B => prdata_13_sqmuxa, 
        C => \addr_data_f0_m_i[6]\, Y => \prdata_39_0_iv_2[6]\);
    
    \reg_sp.addr_matrix_f2[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[4]\);
    
    \reg_wp.delta_f2_f1[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[2]\);
    
    \prdata_RNO_5[10]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[10]\, 
        C => \addr_data_f2_m_i[10]\, Y => \prdata_39_0_iv_3[10]\);
    
    \prdata_RNO_2[10]\ : NOR3C
      port map(A => \prdata_39_0_iv_2[10]\, B => 
        \nb_snapshot_param_m_i[10]\, C => \prdata_39_0_iv_5[10]\, 
        Y => \prdata_39_0_iv_8[10]\);
    
    \prdata_RNO_16[5]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[5]\, 
        Y => \addr_data_f2_m_i[5]\);
    
    \prdata_RNO_3[15]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[15]\, Y => \addr_matrix_f0_1_m_i[15]\);
    
    \apbo.pirq_RNO_3[15]\ : NOR2
      port map(A => status_full_err_0(2), B => 
        status_full_err_0(3), Y => \pirq_2_i_a2_3[15]\);
    
    \prdata_RNO_2[4]\ : NOR3C
      port map(A => \nb_burst_available_m_i[4]\, B => 
        \prdata_39_0_iv_9[4]\, C => data_shaping_R1_m_i, Y => 
        \prdata_39_0_iv_14[4]\);
    
    \prdata_RNO_16[3]\ : OR2B
      port map(A => \status_full_0[3]\, B => prdata_13_sqmuxa, Y
         => \status_full_m_i[3]\);
    
    \prdata_RNO_12[9]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[9]\, 
        Y => \addr_matrix_f2_m_i[9]\);
    
    \reg_sp.addr_matrix_f0_1[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[0]\);
    
    \reg_wp.addr_data_f2[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[0]\);
    
    \reg_wp.addr_data_f2[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[12]\);
    
    \reg_sp.addr_matrix_f1[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[23]\);
    
    \prdata_RNO_4[27]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[27]\, Y
         => \addr_data_f1_m_i[27]\);
    
    \prdata_RNO_0[1]\ : NOR3C
      port map(A => \prdata_39_0_iv_4[1]\, B => 
        \prdata_39_0_iv_3[1]\, C => data_shaping_SP0_m_i, Y => 
        \prdata_39_0_iv_13[1]\);
    
    \prdata[10]\ : DFN1C0
      port map(D => \prdata_39[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(10));
    
    \reg_sp.status_ready_matrix_f1\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_ready_matrix_f1);
    
    \prdata_RNO_0[12]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[12]\, C
         => \addr_data_f1_m_i[12]\, Y => \prdata_39_0_iv_2[12]\);
    
    \prdata_RNO_2[7]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[7]\, B => 
        \prdata_39_0_iv_2[7]\, C => \nb_burst_available_m_i[7]\, 
        Y => \prdata_39_0_iv_10[7]\);
    
    \reg_wp.addr_data_f0[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[4]\);
    
    prdata_2_sqmuxa_0_a2 : NOR3B
      port map(A => N_159, B => N_928, C => apbi_c_19, Y => 
        prdata_2_sqmuxa);
    
    \prdata_RNO[1]\ : OR3C
      port map(A => \prdata_39_0_iv_13[1]\, B => 
        \prdata_39_0_iv_12[1]\, C => \prdata_39_0_iv_14[1]\, Y
         => \prdata_39[1]\);
    
    \prdata_RNO_1[5]\ : AOI1B
      port map(A => \nb_snapshot_param[5]\, B => prdata_18_sqmuxa, 
        C => \prdata_39_0_iv_6[5]\, Y => \prdata_39_0_iv_10[5]\);
    
    \reg_sp.addr_matrix_f0_1[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[28]\);
    
    \reg_sp.addr_matrix_f0_0[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[14]\);
    
    \prdata_RNO_1[2]\ : AOI1B
      port map(A => \nb_burst_available[2]\, B => 
        prdata_17_sqmuxa, C => \prdata_39_0_iv_7[2]\, Y => 
        \prdata_39_0_iv_11[2]\);
    
    \reg_sp.addr_matrix_f0_0[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[15]\);
    
    \reg_sp.addr_matrix_f0_0[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[1]\);
    
    \prdata_RNO_1[24]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[24]\, C
         => \addr_data_f1_m_i[24]\, Y => \prdata_39_0_iv_2[24]\);
    
    \reg_sp.addr_matrix_f0_1[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[30]\);
    
    \reg_sp.addr_matrix_f1_1_sqmuxa_0_a2\ : NOR3B
      port map(A => N_930, B => N_172, C => apbi_c_20, Y => 
        addr_matrix_f1_1_sqmuxa);
    
    \prdata_RNO_0[27]\ : AOI1B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[27]\, C
         => \addr_data_f2_m_i[27]\, Y => \prdata_39_0_iv_3[27]\);
    
    \prdata[13]\ : DFN1C0
      port map(D => \prdata_39[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(13));
    
    \reg_wp.delta_f2_f0[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[3]\);
    
    \reg_wp.enable_f0\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \enable_f0\);
    
    \reg_sp.addr_matrix_f1[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[15]\);
    
    \prdata_RNO_8[15]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[15]\, Y
         => \addr_data_f0_m_i[15]\);
    
    \prdata_RNO_3[18]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[18]\, Y
         => \addr_matrix_f2_m_i[18]\);
    
    \prdata_RNO[15]\ : OR3C
      port map(A => \prdata_39_0_iv_4[15]\, B => 
        \prdata_39_0_iv_3[15]\, C => \prdata_39_0_iv_5[15]\, Y
         => \prdata_39[15]\);
    
    \prdata_RNO_4[10]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[10]\, Y
         => \addr_data_f3_m_i[10]\);
    
    \reg_wp.addr_data_f3[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[0]\);
    
    \prdata_RNO_7[11]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[11]\, Y
         => \addr_data_f0_m_i[11]\);
    
    \reg_wp.addr_data_f0[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[5]\);
    
    \prdata_RNO_7[16]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[16]\, 
        C => \addr_matrix_f2_m_i[16]\, Y => 
        \prdata_39_0_iv_1[16]\);
    
    \reg_sp.addr_matrix_f1[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[12]\);
    
    \prdata[3]\ : DFN1C0
      port map(D => \prdata_39[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(3));
    
    \reg_wp.addr_data_f2[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[27]\);
    
    \reg_wp.burst_f0\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \burst_f0\);
    
    \prdata_RNO_10[4]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[4]\, Y
         => \addr_data_f1_m_i[4]\);
    
    \reg_wp.addr_data_f3[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[15]\);
    
    \prdata[5]\ : DFN1C0
      port map(D => \prdata_39[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(5));
    
    \reg_sp.addr_matrix_f1[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[17]\);
    
    \reg_wp.addr_data_f3[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[16]\);
    
    \prdata_RNO_6[21]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[21]\, Y
         => \addr_data_f2_m_i[21]\);
    
    \prdata_RNO_11[8]\ : OR2B
      port map(A => \nb_burst_available[8]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[8]\);
    
    \prdata_RNO_6[26]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[26]\, 
        Y => \addr_matrix_f0_0_m_i[26]\);
    
    \reg_wp.addr_data_f0[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[24]\);
    
    \prdata_RNO_15[7]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[7]\, Y
         => \delta_f2_f1_m_i[7]\);
    
    \reg_sp.addr_matrix_f2[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[9]\);
    
    \prdata_RNO_7[5]\ : AOI1B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[5]\, C
         => \delta_f2_f1_m_i[5]\, Y => \prdata_39_0_iv_5[5]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \prdata_RNO_2[1]\ : NOR3C
      port map(A => \prdata_39_0_iv_7[1]\, B => 
        \prdata_39_0_iv_6[1]\, C => \prdata_39_0_iv_10[1]\, Y => 
        \prdata_39_0_iv_14[1]\);
    
    \reg_wp.status_new_err[0]\ : DFN1C0
      port map(D => \status_new_err_RNO[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_new_err[0]\);
    
    \reg_wp.status_new_err_RNO[0]\ : OA1B
      port map(A => apbi_c_58, B => \status_full_5_i_o2[0]\, C
         => N_147, Y => \status_new_err_RNO[0]\);
    
    \prdata_RNO_7[12]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[12]\, 
        Y => \addr_matrix_f2_m_i[12]\);
    
    \prdata_RNO_9[2]\ : OR3B
      port map(A => N_161_0, B => \data_shaping_SP1\, C => N_163, 
        Y => data_shaping_SP1_m_i);
    
    \reg_wp.status_full[1]\ : DFN1C0
      port map(D => \status_full_RNO[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \status_full_0[1]\);
    
    \reg_wp.addr_data_f0[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[0]\);
    
    \prdata_RNO_8[18]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[18]\, Y
         => \addr_data_f1_m_i[18]\);
    
    \reg_sp.config_active_interruption_onError_0_sqmuxa_0_o2\ : 
        NOR3A
      port map(A => apbi_c_0, B => apbi_c_24, C => apbi_c_23, Y
         => N_928);
    
    \reg_sp.addr_matrix_f1[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[28]\);
    
    \prdata_RNO_7[8]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[8]\, Y
         => \addr_data_f3_m_i[8]\);
    
    \reg_wp.addr_data_f0[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[28]\);
    
    \prdata_RNO_14[1]\ : OR2B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[1]\, Y
         => \addr_matrix_f1_m_i[1]\);
    
    \reg_wp.delta_snapshot[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[5]\);
    
    \prdata_RNO_2[20]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[20]\, B => 
        \addr_matrix_f0_0_m_i[20]\, C => \prdata_39_0_iv_1[20]\, 
        Y => \prdata_39_0_iv_4[20]\);
    
    \prdata_RNO_6[22]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[22]\, 
        Y => \addr_matrix_f0_0_m_i[22]\);
    
    \prdata_RNO_10[11]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[11]\, 
        Y => \addr_matrix_f2_m_i[11]\);
    
    \reg_wp.nb_snapshot_param[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[0]\);
    
    \prdata_RNO_3[9]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[9]\, Y
         => \delta_snapshot_m_i[9]\);
    
    \reg_wp.addr_data_f0[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[14]\);
    
    \prdata_RNO_1[31]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[31]\, C
         => \addr_data_f1_m_i[31]\, Y => \prdata_39_0_iv_2[31]\);
    
    \prdata_RNO_6[8]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[8]\, Y
         => \delta_f2_f0_m_i[8]\);
    
    \prdata_RNO_5[30]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[30]\, 
        Y => \addr_matrix_f0_1_m_i[30]\);
    
    \prdata_RNO_4[7]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[7]\, 
        C => \addr_matrix_f2_m_i[7]\, Y => \prdata_39_0_iv_1[7]\);
    
    \reg_sp.addr_matrix_f0_1[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[16]\);
    
    \prdata_RNO_5[29]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[29]\, 
        Y => \addr_matrix_f0_1_m_i[29]\);
    
    \prdata_RNO_5[4]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[4]\, C
         => \prdata_39_0_iv_2[4]\, Y => \prdata_39_0_iv_7[4]\);
    
    \prdata_RNO_1[9]\ : NOR3C
      port map(A => \delta_f2_f0_m_i[9]\, B => 
        \addr_data_f3_m_i[9]\, C => \nb_snapshot_param_m_i[9]\, Y
         => \prdata_39_0_iv_8[9]\);
    
    \reg_wp.addr_data_f2[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[1]\);
    
    \reg_wp.delta_f2_f0[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[5]\);
    
    \prdata_RNO_3[17]\ : OR3C
      port map(A => N_161, B => N_168_0, C => \addr_data_f2[17]\, 
        Y => \addr_data_f2_m_i[17]\);
    
    \prdata_RNO_1[23]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[23]\, C => \addr_matrix_f0_1_m_i[23]\, 
        Y => \prdata_39_0_iv_0[23]\);
    
    \prdata_RNO[2]\ : OR3C
      port map(A => \prdata_39_0_iv_12[2]\, B => 
        \prdata_39_0_iv_11[2]\, C => \prdata_39_0_iv_13[2]\, Y
         => \prdata_39[2]\);
    
    \reg_wp.delta_snapshot[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[6]\);
    
    \prdata[15]\ : DFN1C0
      port map(D => \prdata_39[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(15));
    
    \reg_wp.delta_snapshot[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[8]\);
    
    \reg_wp.nb_burst_available[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[6]\);
    
    \reg_wp.status_full_err_RNO[2]\ : OA1B
      port map(A => apbi_c_56, B => \status_full_5_i_o2[0]\, C
         => N_143, Y => \status_full_err_RNO[2]\);
    
    \reg_wp.addr_data_f1[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[23]\);
    
    \reg_wp.addr_data_f0[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[18]\);
    
    \reg_wp.addr_data_f1[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[20]\);
    
    \prdata[6]\ : DFN1C0
      port map(D => \prdata_39[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(6));
    
    \prdata_RNO_4[3]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[3]\, C
         => status_ready_matrix_f2_m_i, Y => 
        \prdata_39_0_iv_2[3]\);
    
    \prdata_RNO_10[9]\ : AOI1B
      port map(A => \status_new_err[1]\, B => prdata_13_sqmuxa, C
         => \addr_data_f0_m_i[9]\, Y => \prdata_39_0_iv_2[9]\);
    
    \reg_wp.status_new_err_RNO[2]\ : OA1B
      port map(A => apbi_c_60, B => \status_full_5_i_o2[0]\, C
         => N_151, Y => \status_new_err_RNO[2]\);
    
    \prdata_RNO_11[6]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[6]\, 
        Y => \addr_matrix_f0_1_m_i[6]\);
    
    \reg_sp.addr_matrix_f0_0[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[22]\);
    
    \reg_wp.status_new_err[2]\ : DFN1C0
      port map(D => \status_new_err_RNO[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_new_err[2]\);
    
    \prdata_RNO_17[4]\ : AOI1B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[4]\, C
         => \delta_f2_f1_m_i[4]\, Y => \prdata_39_0_iv_5[4]\);
    
    \reg_wp.addr_data_f0[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[3]\);
    
    \reg_wp.addr_data_f3[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[12]\);
    
    \prdata_RNO_0[6]\ : AOI1B
      port map(A => \nb_burst_available[6]\, B => 
        prdata_17_sqmuxa, C => \prdata_39_0_iv_6[6]\, Y => 
        \prdata_39_0_iv_10[6]\);
    
    prdata_4_sqmuxa_0_a2_0 : NOR2B
      port map(A => N_172, B => N_161_0, Y => prdata_4_sqmuxa_0);
    
    \reg_wp.delta_f2_f1[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[3]\);
    
    \prdata_RNO_8[24]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[24]\, Y
         => \addr_matrix_f2_m_i[24]\);
    
    \reg_wp.addr_data_f1[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[21]\);
    
    \prdata_RNO_2[0]\ : NOR3C
      port map(A => \prdata_39_0_iv_4[0]\, B => 
        \prdata_39_0_iv_3[0]\, C => \prdata_39_0_iv_11[0]\, Y => 
        \prdata_39_0_iv_14[0]\);
    
    \reg_wp.delta_f2_f0[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[8]\);
    
    \reg_wp.addr_data_f2[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[9]\);
    
    \prdata_RNO[27]\ : OR3C
      port map(A => \prdata_39_0_iv_3[27]\, B => 
        \prdata_39_0_iv_2[27]\, C => \prdata_39_0_iv_4[27]\, Y
         => \prdata_39[27]\);
    
    \prdata_RNO_8[30]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[30]\, Y
         => \addr_matrix_f2_m_i[30]\);
    
    \prdata_RNO_3[29]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[29]\, Y
         => \addr_data_f2_m_i[29]\);
    
    prdata_4_sqmuxa_0_a2 : NOR2B
      port map(A => N_172, B => N_161, Y => prdata_4_sqmuxa);
    
    \prdata_RNO_8[17]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[17]\, Y
         => \addr_matrix_f2_m_i[17]\);
    
    \reg_wp.status_full_RNO_0[3]\ : NOR3A
      port map(A => N_933_0, B => \status_full_0[3]\, C => 
        status_full(3), Y => N_138);
    
    \prdata_RNO_18[2]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[2]\, 
        C => \addr_matrix_f2_m_i[2]\, Y => \prdata_39_0_iv_1[2]\);
    
    \apbo.pirq_RNO_1[15]\ : NOR3A
      port map(A => \pirq_2_i_a2_1[15]\, B => status_new_err_0_1, 
        C => status_new_err_0_0, Y => \pirq_2_i_a2_6[15]\);
    
    \reg_wp.status_full_err_RNO_0[0]\ : NOR3A
      port map(A => N_933_0, B => \status_full_err[0]\, C => 
        status_full_err_0(0), Y => N_139);
    
    \prdata_RNO_6[14]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[14]\, 
        C => \addr_data_f2_m_i[14]\, Y => \prdata_39_0_iv_3[14]\);
    
    \prdata_RNO_1[11]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[11]\, B => 
        \addr_matrix_f0_0_m_i[11]\, C => \addr_data_f3_m_i[11]\, 
        Y => \prdata_39_0_iv_4[11]\);
    
    \prdata_RNO_1[16]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[16]\, C
         => \addr_data_f1_m_i[16]\, Y => \prdata_39_0_iv_2[16]\);
    
    \apbo.pirq[15]\ : DFN1C0
      port map(D => N_155_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => pirq_c(15));
    
    \reg_wp.addr_data_f1[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[4]\);
    
    \prdata_RNO[19]\ : OR3C
      port map(A => \prdata_39_0_iv_3[19]\, B => 
        \prdata_39_0_iv_2[19]\, C => \prdata_39_0_iv_4[19]\, Y
         => \prdata_39[19]\);
    
    \reg_wp.data_shaping_BW\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => \data_shaping_BW_c\);
    
    \reg_wp.delta_f2_f0_1_sqmuxa_0_a2_0\ : NOR3A
      port map(A => N_158, B => apbi_c_21, C => apbi_c_22, Y => 
        N_164);
    
    \prdata_RNO_17[1]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[1]\, 
        Y => \addr_matrix_f0_0_m_i[1]\);
    
    \reg_sp.addr_matrix_f2[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[0]\);
    
    \prdata_RNO_9[1]\ : AOI1B
      port map(A => \nb_snapshot_param[1]\, B => prdata_18_sqmuxa, 
        C => \prdata_39_0_iv_5[1]\, Y => \prdata_39_0_iv_10[1]\);
    
    \prdata_RNO_1[0]\ : AOI1B
      port map(A => \nb_snapshot_param[0]\, B => prdata_18_sqmuxa, 
        C => \prdata_39_0_iv_7[0]\, Y => \prdata_39_0_iv_12[0]\);
    
    \prdata_RNO_10[1]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[1]\, 
        Y => \addr_data_f2_m_i[1]\);
    
    \reg_sp.addr_matrix_f0_0_1_sqmuxa_0_a2_0\ : NOR3C
      port map(A => N_159, B => N_928, C => N_930, Y => 
        addr_matrix_f0_0_1_sqmuxa_0);
    
    \reg_wp.addr_data_f1[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[13]\);
    
    \reg_wp.delta_snapshot[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[4]\);
    
    \reg_wp.addr_data_f1[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[10]\);
    
    \reg_wp.status_full_RNO_0[0]\ : NOR3A
      port map(A => N_933_0, B => \status_full_0[0]\, C => 
        status_full(0), Y => N_135);
    
    \reg_sp.addr_matrix_f1[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[9]\);
    
    \reg_wp.delta_f2_f1[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[8]\);
    
    \reg_sp.addr_matrix_f0_1[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[10]\);
    
    \prdata_RNO_19[3]\ : OR2B
      port map(A => \nb_burst_available[3]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[3]\);
    
    \prdata_RNO_2[5]\ : NOR3C
      port map(A => \prdata_39_0_iv_5[5]\, B => 
        \prdata_39_0_iv_4[5]\, C => \nb_burst_available_m_i[5]\, 
        Y => \prdata_39_0_iv_12[5]\);
    
    \prdata_RNO_2[6]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[6]\, B => 
        \prdata_39_0_iv_2[6]\, C => \prdata_39_0_iv_8[6]\, Y => 
        \prdata_39_0_iv_11[6]\);
    
    prdata_8_sqmuxa_0_a2 : NOR2
      port map(A => N_163, B => N_157, Y => prdata_8_sqmuxa);
    
    \prdata_RNO_0[19]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[19]\, 
        C => \addr_data_f2_m_i[19]\, Y => \prdata_39_0_iv_3[19]\);
    
    \prdata[12]\ : DFN1C0
      port map(D => \prdata_39[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(12));
    
    \reg_sp.addr_matrix_f0_1[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[13]\);
    
    \prdata_RNO_1[12]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[12]\, 
        Y => \delta_snapshot_m_i[12]\);
    
    \reg_sp.addr_matrix_f0_0[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[9]\);
    
    \reg_wp.addr_data_f1[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[11]\);
    
    prdata_0_sqmuxa_0_a2 : NOR2A
      port map(A => N_161, B => N_169, Y => prdata_0_sqmuxa);
    
    \prdata_RNO_5[25]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[25]\, 
        Y => \addr_matrix_f0_1_m_i[25]\);
    
    \prdata[19]\ : DFN1C0
      port map(D => \prdata_39[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(19));
    
    \prdata_RNO_11[4]\ : AOI1B
      port map(A => \status_full_err[0]\, B => prdata_13_sqmuxa, 
        C => status_error_anticipating_empty_fifo_m_i, Y => 
        \prdata_39_0_iv_2[4]\);
    
    \reg_wp.delta_f2_f0[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[7]\);
    
    \prdata_RNO_11[11]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[11]\, Y => \addr_data_f2_m_i[11]\);
    
    \reg_sp.addr_matrix_f0_1[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[29]\);
    
    \reg_wp.status_full_RNO[1]\ : OA1B
      port map(A => apbi_c_51, B => \status_full_5_i_o2[0]\, C
         => N_136, Y => \status_full_RNO[1]\);
    
    \reg_wp.nb_burst_available[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[5]\);
    
    \prdata_RNO_7[30]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[30]\, C
         => \addr_matrix_f2_m_i[30]\, Y => \prdata_39_0_iv_1[30]\);
    
    \reg_wp.addr_data_f3[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[8]\);
    
    \prdata_RNO_5[11]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[11]\, 
        Y => \addr_matrix_f0_0_m_i[11]\);
    
    \reg_wp.addr_data_f0[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[29]\);
    
    \prdata_RNO_5[16]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[16]\, Y => \addr_matrix_f0_1_m_i[16]\);
    
    \prdata_RNO_2[11]\ : NOR3C
      port map(A => \addr_data_f0_m_i[11]\, B => 
        \status_new_err_m_i[3]\, C => \prdata_39_0_iv_3[11]\, Y
         => \prdata_39_0_iv_6[11]\);
    
    \prdata_RNO_2[16]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[16]\, B => 
        \addr_matrix_f0_0_m_i[16]\, C => \prdata_39_0_iv_1[16]\, 
        Y => \prdata_39_0_iv_4[16]\);
    
    \prdata_RNO_13[10]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[10]\, 
        Y => \addr_matrix_f2_m_i[10]\);
    
    \reg_wp.nb_burst_available[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[8]\);
    
    \reg_wp.addr_data_f2_1_sqmuxa_0_a2\ : NOR3B
      port map(A => N_930, B => N_168, C => apbi_c_20, Y => 
        addr_data_f2_1_sqmuxa);
    
    prdata_13_sqmuxa_0_a2 : NOR3A
      port map(A => apbi_c_21, B => N_931, C => apbi_c_19, Y => 
        prdata_13_sqmuxa);
    
    \reg_wp.delta_f2_f0[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[0]\);
    
    \reg_sp.status_error_bad_component_error\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_error_bad_component_error);
    
    \prdata_RNO_12[10]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[10]\, 
        C => \addr_matrix_f2_m_i[10]\, Y => 
        \prdata_39_0_iv_1[10]\);
    
    \reg_wp.addr_data_f3[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[24]\);
    
    \reg_wp.nb_burst_available[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[4]\);
    
    prdata_10_sqmuxa_0_a2_0 : NOR3A
      port map(A => apbi_c_19, B => apbi_c_21, C => N_931, Y => 
        prdata_10_sqmuxa_0);
    
    \reg_wp.addr_data_f1[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[25]\);
    
    \lpp_top_apbreg.reg_wp.status_full_5_i_o2_0[0]\ : OR3B
      port map(A => apbi_c_21, B => N_930, C => N_931, Y => 
        N_933_0);
    
    \reg_wp.addr_data_f1[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[26]\);
    
    \prdata_RNO_0[30]\ : AOI1B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[30]\, C
         => \addr_data_f2_m_i[30]\, Y => \prdata_39_0_iv_3[30]\);
    
    \reg_wp.addr_data_f1[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[1]\);
    
    \prdata_RNO_8[23]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[23]\, Y
         => \addr_data_f1_m_i[23]\);
    
    \reg_sp.addr_matrix_f2[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[3]\);
    
    \reg_sp.addr_matrix_f2[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[19]\);
    
    \status_full_ack[0]\ : DFN1C0
      port map(D => \status_full_ack_8[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => status_full_ack(0));
    
    \prdata[21]\ : DFN1C0
      port map(D => \prdata_39[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(21));
    
    \prdata_RNO_3[8]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[8]\, 
        C => \addr_matrix_f0_1_m_i[8]\, Y => 
        \prdata_39_0_iv_0[8]\);
    
    \prdata_RNO_5[12]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[12]\, C => \addr_matrix_f0_1_m_i[12]\, 
        Y => \prdata_39_0_iv_0[12]\);
    
    \reg_wp.addr_data_f3[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[28]\);
    
    \reg_wp.addr_data_f2[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[23]\);
    
    \prdata_RNO_5[28]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[28]\, 
        Y => \addr_matrix_f0_1_m_i[28]\);
    
    \prdata_RNO_2[12]\ : NOR3C
      port map(A => \prdata_39_0_iv_1[12]\, B => 
        \prdata_39_0_iv_0[12]\, C => \prdata_39_0_iv_3[12]\, Y
         => \prdata_39_0_iv_6[12]\);
    
    \reg_wp.addr_data_f2[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[20]\);
    
    \prdata_RNO_1[20]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[20]\, C
         => \addr_data_f1_m_i[20]\, Y => \prdata_39_0_iv_2[20]\);
    
    \prdata_RNO_10[0]\ : OR3A
      port map(A => status_ready_matrix_f0_0, B => N_157, C => 
        N_169, Y => status_ready_matrix_f0_0_m_i);
    
    \reg_wp.data_shaping_SP0\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => \data_shaping_SP0\);
    
    \prdata_RNO_6[13]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[13]\, 
        C => \addr_data_f2_m_i[13]\, Y => \prdata_39_0_iv_3[13]\);
    
    \prdata_RNO_3[25]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[25]\, Y
         => \addr_data_f2_m_i[25]\);
    
    \reg_wp.addr_data_f0[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[19]\);
    
    \prdata_RNO_11[9]\ : OR2B
      port map(A => \nb_burst_available[9]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[9]\);
    
    \prdata_RNO_17[9]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[9]\, Y
         => \addr_data_f0_m_i[9]\);
    
    \reg_wp.data_shaping_R1_0\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => \data_shaping_R1_0\);
    
    \prdata_RNO_8[5]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[5]\, C
         => \addr_data_f2_m_i[5]\, Y => \prdata_39_0_iv_4[5]\);
    
    \prdata_RNO_6[3]\ : OR2B
      port map(A => \nb_snapshot_param[3]\, B => prdata_18_sqmuxa, 
        Y => \nb_snapshot_param_m_i[3]\);
    
    \reg_sp.addr_matrix_f2[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[13]\);
    
    \prdata_RNO_17[6]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[6]\, Y
         => \addr_data_f3_m_i[6]\);
    
    \prdata_RNO_7[19]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[19]\, C
         => \addr_matrix_f2_m_i[19]\, Y => \prdata_39_0_iv_1[19]\);
    
    \prdata_RNO_9[14]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[14]\, Y
         => \addr_data_f2_m_i[14]\);
    
    \prdata_RNO_7[24]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[24]\, C
         => \addr_matrix_f2_m_i[24]\, Y => \prdata_39_0_iv_1[24]\);
    
    \prdata_RNO[21]\ : OR3C
      port map(A => \prdata_39_0_iv_1[21]\, B => 
        \prdata_39_0_iv_0[21]\, C => \prdata_39_0_iv_5[21]\, Y
         => \prdata_39[21]\);
    
    \prdata[1]\ : DFN1C0
      port map(D => \prdata_39[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(1));
    
    \reg_wp.delta_snapshot[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[10]\);
    
    \reg_sp.addr_matrix_f2[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[29]\);
    
    \reg_wp.addr_data_f2[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[21]\);
    
    \reg_wp.addr_data_f3[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[7]\);
    
    \prdata_RNO_4[11]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[11]\, Y => \addr_matrix_f0_1_m_i[11]\);
    
    \prdata_RNO_4[16]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[16]\, 
        Y => \addr_data_f1_m_i[16]\);
    
    \prdata_RNO_1[7]\ : NOR3C
      port map(A => \delta_f2_f0_m_i[7]\, B => 
        \addr_data_f3_m_i[7]\, C => \nb_snapshot_param_m_i[7]\, Y
         => \prdata_39_0_iv_8[7]\);
    
    \prdata_RNO_7[9]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[9]\, Y
         => \addr_data_f3_m_i[9]\);
    
    \prdata_RNO_6[29]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[29]\, 
        Y => \addr_matrix_f0_0_m_i[29]\);
    
    \prdata_RNO_19[2]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[2]\, Y
         => \delta_f2_f0_m_i[2]\);
    
    \reg_wp.addr_data_f1[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[15]\);
    
    \prdata_RNO_16[2]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[2]\, 
        Y => \addr_matrix_f0_1_m_i[2]\);
    
    \reg_wp.status_full_err_RNO[0]\ : OA1B
      port map(A => apbi_c_54, B => \status_full_5_i_o2[0]\, C
         => N_139, Y => \status_full_err_RNO[0]\);
    
    \reg_wp.addr_data_f1[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[16]\);
    
    \prdata_RNO_5[9]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[9]\, B => 
        \addr_matrix_f0_0_m_i[9]\, C => \delta_f2_f1_m_i[9]\, Y
         => \prdata_39_0_iv_5[9]\);
    
    \reg_sp.addr_matrix_f1[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[26]\);
    
    \reg_sp.addr_matrix_f2[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[2]\);
    
    \reg_sp.addr_matrix_f0_1[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[14]\);
    
    \reg_sp.addr_matrix_f0_1[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[15]\);
    
    \prdata_RNO[26]\ : OR3C
      port map(A => \prdata_39_0_iv_3[26]\, B => 
        \prdata_39_0_iv_2[26]\, C => \prdata_39_0_iv_4[26]\, Y
         => \prdata_39[26]\);
    
    \prdata_RNO_0[15]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[15]\, B => 
        \addr_matrix_f0_0_m_i[15]\, C => \prdata_39_0_iv_1[15]\, 
        Y => \prdata_39_0_iv_4[15]\);
    
    \prdata[31]\ : DFN1C0
      port map(D => \prdata_39[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(31));
    
    \reg_wp.addr_data_f1_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_166, B => apbi_c_21, C => N_931, Y => 
        addr_data_f1_1_sqmuxa);
    
    \reg_wp.addr_data_f2[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[30]\);
    
    \reg_sp.addr_matrix_f0_1[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[7]\);
    
    \prdata_RNO_4[24]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[24]\, Y
         => \addr_data_f1_m_i[24]\);
    
    \reg_sp.addr_matrix_f1[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[21]\);
    
    \reg_sp.addr_matrix_f2[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[23]\);
    
    \reg_wp.addr_data_f3[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[3]\);
    
    \prdata_RNO_3[28]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[28]\, Y
         => \addr_data_f2_m_i[28]\);
    
    \reg_sp.addr_matrix_f1[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[20]\);
    
    \prdata[16]\ : DFN1C0
      port map(D => \prdata_39[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(16));
    
    \prdata_RNO_4[0]\ : AOI1B
      port map(A => prdata_0_sqmuxa, B => 
        config_active_interruption_onNewMatrix, C => 
        status_ready_matrix_f0_0_m_i, Y => \prdata_39_0_iv_2[0]\);
    
    \status_full_ack[2]\ : DFN1C0
      port map(D => \status_full_ack_8[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => status_full_ack(2));
    
    \prdata_RNO_4[12]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[12]\, 
        C => \addr_matrix_f2_m_i[12]\, Y => 
        \prdata_39_0_iv_1[12]\);
    
    \prdata_RNO[0]\ : OR3C
      port map(A => \prdata_39_0_iv_13[0]\, B => 
        \prdata_39_0_iv_12[0]\, C => \prdata_39_0_iv_14[0]\, Y
         => \prdata_39[0]\);
    
    \reg_wp.addr_data_f1[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[22]\);
    
    \prdata_RNO_12[5]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[5]\, 
        Y => \addr_matrix_f0_1_m_i[5]\);
    
    \reg_wp.addr_data_f2[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[31]\);
    
    \reg_wp.nb_snapshot_param[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[3]\);
    
    \reg_sp.addr_matrix_f0_0[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[12]\);
    
    \prdata_RNO_0[24]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[24]\, 
        C => \addr_data_f2_m_i[24]\, Y => \prdata_39_0_iv_3[24]\);
    
    \reg_sp.status_error_anticipating_empty_fifo\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_error_anticipating_empty_fifo);
    
    \reg_sp.addr_matrix_f0_0[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[8]\);
    
    \status_full_ack_RNO[0]\ : NOR3A
      port map(A => \status_full_0[0]\, B => apbi_c_50, C => 
        \status_full_5_i_o2[0]\, Y => \status_full_ack_8[0]\);
    
    \prdata_RNO_2[21]\ : NOR3C
      port map(A => \addr_data_f3_m_i[21]\, B => 
        \addr_data_f2_m_i[21]\, C => \prdata_39_0_iv_2[21]\, Y
         => \prdata_39_0_iv_5[21]\);
    
    \reg_sp.addr_matrix_f0_0[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[21]\);
    
    \prdata_RNO_2[26]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[26]\, B => 
        \addr_matrix_f0_0_m_i[26]\, C => \prdata_39_0_iv_1[26]\, 
        Y => \prdata_39_0_iv_4[26]\);
    
    \prdata_RNO_5[27]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[27]\, 
        Y => \addr_matrix_f0_1_m_i[27]\);
    
    \reg_wp.addr_data_f0[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[2]\);
    
    \reg_sp.addr_matrix_f0_0[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[0]\);
    
    \prdata_RNO_5[1]\ : OR3B
      port map(A => N_161_0, B => \data_shaping_SP0\, C => N_163, 
        Y => data_shaping_SP0_m_i);
    
    \prdata_RNO_15[8]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[8]\, Y
         => \delta_snapshot_m_i[8]\);
    
    \prdata_RNO_15[6]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[6]\, Y
         => \addr_data_f0_m_i[6]\);
    
    \reg_wp.status_full[3]\ : DFN1C0
      port map(D => \status_full_RNO[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \status_full_0[3]\);
    
    \prdata_RNO_16[1]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[1]\, 
        Y => \addr_matrix_f0_1_m_i[1]\);
    
    \prdata[2]\ : DFN1C0
      port map(D => \prdata_39[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(2));
    
    \reg_wp.delta_snapshot[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[2]\);
    
    \prdata_RNO_5[31]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[31]\, 
        Y => \addr_matrix_f0_1_m_i[31]\);
    
    prdata_9_sqmuxa_0_a2 : NOR3
      port map(A => apbi_c_21, B => N_931, C => apbi_c_19, Y => 
        prdata_9_sqmuxa);
    
    \prdata_RNO_5[2]\ : NOR3C
      port map(A => \status_full_m_i[2]\, B => 
        \delta_f2_f1_m_i[2]\, C => \prdata_39_0_iv_4[2]\, Y => 
        \prdata_39_0_iv_9[2]\);
    
    \prdata_RNO_0[18]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[18]\, 
        C => \addr_matrix_f2_m_i[18]\, Y => 
        \prdata_39_0_iv_1[18]\);
    
    \reg_wp.nb_snapshot_param[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[6]\);
    
    \reg_wp.addr_data_f2_1_sqmuxa_0_a2_0_1\ : NOR3B
      port map(A => N_930, B => N_168, C => apbi_c_20, Y => 
        addr_data_f2_1_sqmuxa_0);
    
    \reg_sp.addr_matrix_f2[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[18]\);
    
    \lpp_top_apbreg.reg_wp.status_full_5_i_o2[0]\ : OR3B
      port map(A => apbi_c_21, B => N_930, C => N_931, Y => 
        \status_full_5_i_o2[0]\);
    
    \reg_wp.status_new_err_RNO_0[0]\ : NOR3A
      port map(A => N_933_0, B => \status_new_err[0]\, C => 
        status_new_err_0_0, Y => N_147);
    
    \reg_wp.delta_f2_f1[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[6]\);
    
    \reg_sp.addr_matrix_f0_1[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[27]\);
    
    \reg_wp.status_full_err[0]\ : DFN1C0
      port map(D => \status_full_err_RNO[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_full_err[0]\);
    
    \prdata_RNO_18[3]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[3]\, 
        C => \addr_matrix_f2_m_i[3]\, Y => \prdata_39_0_iv_1[3]\);
    
    \reg_sp.addr_matrix_f1[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[4]\);
    
    \reg_sp.addr_matrix_f1[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[19]\);
    
    \reg_wp.addr_data_f2[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[25]\);
    
    \prdata_RNO_9[9]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[9]\, C
         => \addr_data_f2_m_i[9]\, Y => \prdata_39_0_iv_3[9]\);
    
    \prdata_RNO_9[13]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[13]\, Y => \addr_data_f2_m_i[13]\);
    
    \prdata_RNO_3[5]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[5]\, C
         => \addr_data_f1_m_i[5]\, Y => \prdata_39_0_iv_3[5]\);
    
    \prdata_RNO_0[4]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[4]\, B => burst_f0_m_i, C
         => \prdata_39_0_iv_7[4]\, Y => \prdata_39_0_iv_11[4]\);
    
    \prdata_RNO_7[23]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[23]\, C
         => \addr_data_f1_m_i[23]\, Y => \prdata_39_0_iv_2[23]\);
    
    \reg_wp.addr_data_f2[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[26]\);
    
    \prdata_RNO_2[22]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[22]\, B => 
        \addr_matrix_f0_0_m_i[22]\, C => \prdata_39_0_iv_1[22]\, 
        Y => \prdata_39_0_iv_4[22]\);
    
    \reg_sp.addr_matrix_f0_1[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[8]\);
    
    \reg_wp.delta_snapshot[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[7]\);
    
    \reg_sp.addr_matrix_f0_0[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[3]\);
    
    \prdata_RNO_18[6]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \burst_f2\, Y => 
        burst_f2_m_i);
    
    \reg_wp.burst_f1\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \burst_f1\);
    
    \prdata_RNO_7[15]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[15]\, 
        Y => \addr_data_f1_m_i[15]\);
    
    \reg_wp.addr_data_f1[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[12]\);
    
    \reg_sp.addr_matrix_f1[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[7]\);
    
    \reg_wp.status_full_RNO[2]\ : OA1B
      port map(A => apbi_c_52, B => \status_full_5_i_o2[0]\, C
         => N_137, Y => \status_full_RNO[2]\);
    
    \reg_wp.nb_burst_available[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[1]\);
    
    \prdata_RNO_8[20]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[20]\, Y
         => \addr_matrix_f2_m_i[20]\);
    
    \prdata_RNO_0[5]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[5]\, B => burst_f1_m_i, C
         => \prdata_39_0_iv_7[5]\, Y => \prdata_39_0_iv_11[5]\);
    
    \reg_wp.addr_data_f2[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[14]\);
    
    \reg_sp.addr_matrix_f0_0[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[28]\);
    
    \reg_wp.addr_data_f3[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[30]\);
    
    \prdata_RNO_3[27]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[27]\, Y
         => \addr_data_f2_m_i[27]\);
    
    \reg_wp.addr_data_f0[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[1]\);
    
    \reg_sp.addr_matrix_f1[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[13]\);
    
    \prdata_RNO_6[25]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[25]\, 
        Y => \addr_matrix_f0_0_m_i[25]\);
    
    \reg_wp.addr_data_f3[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[29]\);
    
    \reg_sp.addr_matrix_f2[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[28]\);
    
    \prdata_RNO_12[8]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[8]\, 
        Y => \addr_matrix_f0_1_m_i[8]\);
    
    \prdata_RNO_4[23]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[23]\, 
        Y => \addr_matrix_f0_1_m_i[23]\);
    
    \prdata_RNO_1[19]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[19]\, C
         => \addr_data_f1_m_i[19]\, Y => \prdata_39_0_iv_2[19]\);
    
    \prdata_RNO_8[31]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[31]\, Y
         => \addr_matrix_f2_m_i[31]\);
    
    \prdata_RNO_7[2]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[2]\, B => 
        \addr_matrix_f0_0_m_i[2]\, C => \prdata_39_0_iv_1[2]\, Y
         => \prdata_39_0_iv_6[2]\);
    
    \prdata_RNO_6[10]\ : AOI1B
      port map(A => \status_new_err[2]\, B => prdata_13_sqmuxa, C
         => \addr_data_f0_m_i[10]\, Y => \prdata_39_0_iv_2[10]\);
    
    \reg_sp.addr_matrix_f1[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[24]\);
    
    \prdata_RNO_7[6]\ : NOR3C
      port map(A => \delta_f2_f0_m_i[6]\, B => 
        \addr_data_f3_m_i[6]\, C => burst_f2_m_i, Y => 
        \prdata_39_0_iv_8[6]\);
    
    \reg_wp.data_shaping_BW_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_930, B => apbi_c_20, C => N_163, Y => 
        data_shaping_BW_1_sqmuxa);
    
    \reg_wp.addr_data_f3[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[31]\);
    
    \reg_wp.addr_data_f2[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[18]\);
    
    \prdata_RNO[5]\ : OR3C
      port map(A => \prdata_39_0_iv_11[5]\, B => 
        \prdata_39_0_iv_10[5]\, C => \prdata_39_0_iv_12[5]\, Y
         => \prdata_39[5]\);
    
    \prdata_RNO_3[14]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[14]\, Y
         => \addr_data_f1_m_i[14]\);
    
    \reg_wp.status_full[2]\ : DFN1C0
      port map(D => \status_full_RNO[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \status_full_0[2]\);
    
    \prdata_RNO_0[23]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[23]\, C
         => \addr_matrix_f2_m_i[23]\, Y => \prdata_39_0_iv_1[23]\);
    
    \reg_wp.status_full_RNO[0]\ : OA1B
      port map(A => apbi_c_50, B => \status_full_5_i_o2[0]\, C
         => N_135, Y => \status_full_RNO[0]\);
    
    \prdata_RNO_7[18]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[18]\, C
         => \addr_data_f1_m_i[18]\, Y => \prdata_39_0_iv_2[18]\);
    
    \prdata_RNO_13[9]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[9]\, 
        Y => \addr_matrix_f0_1_m_i[9]\);
    
    \reg_wp.addr_data_f1[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[2]\);
    
    \reg_sp.addr_matrix_f2[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[6]\);
    
    \prdata_RNO_0[17]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[17]\, 
        C => \addr_data_f2_m_i[17]\, Y => \prdata_39_0_iv_3[17]\);
    
    prdata_0_sqmuxa_0_a2_0_0 : NOR2
      port map(A => apbi_c_20, B => apbi_c_19, Y => N_161_0);
    
    \reg_wp.addr_data_f1[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[3]\);
    
    \prdata_RNO_0[9]\ : NOR3C
      port map(A => \delta_snapshot_m_i[9]\, B => 
        \prdata_39_0_iv_1[9]\, C => \prdata_39_0_iv_5[9]\, Y => 
        \prdata_39_0_iv_9[9]\);
    
    \reg_sp.addr_matrix_f0_0[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[30]\);
    
    \prdata_RNO_6[28]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[28]\, 
        Y => \addr_matrix_f0_0_m_i[28]\);
    
    \reg_wp.addr_data_f2[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[3]\);
    
    \prdata_RNO[31]\ : OR3C
      port map(A => \prdata_39_0_iv_3[31]\, B => 
        \prdata_39_0_iv_2[31]\, C => \prdata_39_0_iv_4[31]\, Y
         => \prdata_39[31]\);
    
    \reg_sp.addr_matrix_f0_0[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[6]\);
    
    \prdata_RNO_17[5]\ : OR3A
      port map(A => status_error_bad_component_error, B => N_157, 
        C => N_169, Y => status_error_bad_component_error_m_i);
    
    \prdata_RNO_10[7]\ : AOI1B
      port map(A => \status_full_err[3]\, B => prdata_13_sqmuxa, 
        C => \addr_data_f0_m_i[7]\, Y => \prdata_39_0_iv_2[7]\);
    
    \prdata_RNO_13[4]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[4]\, 
        Y => \addr_matrix_f0_0_m_i[4]\);
    
    \reg_sp.addr_matrix_f1_1_sqmuxa_0_a2_0\ : NOR3B
      port map(A => N_930, B => N_172, C => apbi_c_20, Y => 
        addr_matrix_f1_1_sqmuxa_0);
    
    \reg_sp.addr_matrix_f0_1_1_sqmuxa_0_a2\ : NOR3C
      port map(A => N_159, B => N_928, C => N_166, Y => 
        addr_matrix_f0_1_1_sqmuxa);
    
    \prdata_RNO_5[19]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[19]\, 
        Y => \addr_matrix_f0_1_m_i[19]\);
    
    \prdata_RNO_2[19]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[19]\, B => 
        \addr_matrix_f0_0_m_i[19]\, C => \prdata_39_0_iv_1[19]\, 
        Y => \prdata_39_0_iv_4[19]\);
    
    \prdata_RNO_3[2]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[2]\, C
         => \addr_data_f2_m_i[2]\, Y => \prdata_39_0_iv_3[2]\);
    
    \prdata_RNO_0[7]\ : NOR3C
      port map(A => \delta_snapshot_m_i[7]\, B => 
        \prdata_39_0_iv_1[7]\, C => \prdata_39_0_iv_5[7]\, Y => 
        \prdata_39_0_iv_9[7]\);
    
    \reg_wp.addr_data_f2[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[22]\);
    
    \reg_wp.delta_f2_f0[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[9]\);
    
    \prdata[17]\ : DFN1C0
      port map(D => \prdata_39[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(17));
    
    \reg_wp.addr_data_f0[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[30]\);
    
    \prdata_RNO_7[31]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[31]\, C
         => \addr_matrix_f2_m_i[31]\, Y => \prdata_39_0_iv_1[31]\);
    
    \prdata_RNO_8[2]\ : OR2B
      port map(A => \nb_snapshot_param[2]\, B => prdata_18_sqmuxa, 
        Y => \nb_snapshot_param_m_i[2]\);
    
    \reg_wp.status_full_err[2]\ : DFN1C0
      port map(D => \status_full_err_RNO[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_full_err[2]\);
    
    \prdata_RNO_11[2]\ : OR3A
      port map(A => status_ready_matrix_f1, B => N_157, C => 
        N_169, Y => status_ready_matrix_f1_m_i);
    
    \prdata_RNO_8[14]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[14]\, Y => \addr_matrix_f0_1_m_i[14]\);
    
    \reg_sp.addr_matrix_f2[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[31]\);
    
    \prdata_RNO_15[2]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \enable_f2\, Y => 
        enable_f2_m_i);
    
    \prdata[18]\ : DFN1C0
      port map(D => \prdata_39[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(18));
    
    \reg_sp.addr_matrix_f2[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[30]\);
    
    \reg_wp.addr_data_f2[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[7]\);
    
    \prdata_RNO[13]\ : OR3C
      port map(A => \prdata_39_0_iv_2[13]\, B => 
        \delta_snapshot_m_i[13]\, C => \prdata_39_0_iv_6[13]\, Y
         => \prdata_39[13]\);
    
    \reg_wp.data_shaping_R0_0\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => \data_shaping_R0_0\);
    
    \reg_sp.addr_matrix_f1[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[2]\);
    
    \reg_sp.addr_matrix_f1[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[18]\);
    
    \prdata_RNO_9[3]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[3]\, 
        Y => \addr_data_f2_m_i[3]\);
    
    \prdata_RNO_21[0]\ : OR3B
      port map(A => N_161, B => \data_shaping_BW_c\, C => N_163, 
        Y => data_shaping_BW_m_i);
    
    \prdata_RNO_15[9]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[9]\, Y
         => \delta_f2_f1_m_i[9]\);
    
    \prdata_RNO_0[31]\ : AOI1B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[31]\, C
         => \addr_data_f2_m_i[31]\, Y => \prdata_39_0_iv_3[31]\);
    
    \prdata_RNO_0[3]\ : OR3B
      port map(A => N_161_0, B => \data_shaping_R0_0\, C => N_163, 
        Y => data_shaping_R0_m_i);
    
    \prdata_RNO[3]\ : OR3C
      port map(A => data_shaping_R0_m_i, B => 
        \prdata_39_0_iv_12[3]\, C => \prdata_39_0_iv_13[3]\, Y
         => \prdata_39[3]\);
    
    \reg_wp.enable_f2\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \enable_f2\);
    
    \reg_wp.addr_data_f0[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[6]\);
    
    \reg_wp.addr_data_f0[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[31]\);
    
    \prdata_RNO[6]\ : OR3C
      port map(A => \prdata_39_0_iv_10[6]\, B => 
        \prdata_39_0_iv_9[6]\, C => \prdata_39_0_iv_11[6]\, Y => 
        \prdata_39[6]\);
    
    \reg_wp.status_new_err_RNO_0[1]\ : NOR3A
      port map(A => N_933_0, B => \status_new_err[1]\, C => 
        status_new_err_0_1, Y => N_149);
    
    \reg_wp.addr_data_f3[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[9]\);
    
    \reg_wp.status_new_err[1]\ : DFN1C0
      port map(D => \status_new_err_RNO[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_new_err[1]\);
    
    \prdata_RNO_10[5]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[5]\, Y
         => \addr_data_f1_m_i[5]\);
    
    \prdata_RNO_16[7]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[7]\, 
        Y => \addr_data_f2_m_i[7]\);
    
    \prdata_RNO_1[1]\ : AOI1B
      port map(A => \nb_burst_available[1]\, B => 
        prdata_17_sqmuxa, C => \prdata_39_0_iv_8[1]\, Y => 
        \prdata_39_0_iv_12[1]\);
    
    \reg_wp.status_full_RNO_0[1]\ : NOR3A
      port map(A => N_933_0, B => \status_full_0[1]\, C => 
        status_full(1), Y => N_136);
    
    \prdata_RNO_14[6]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[6]\, 
        Y => \addr_data_f2_m_i[6]\);
    
    \prdata_RNO_1[21]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[21]\, C => \addr_matrix_f0_1_m_i[21]\, 
        Y => \prdata_39_0_iv_0[21]\);
    
    \prdata_RNO_1[26]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[26]\, C
         => \addr_data_f1_m_i[26]\, Y => \prdata_39_0_iv_2[26]\);
    
    \prdata_RNO_1[15]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[15]\, 
        C => \addr_data_f2_m_i[15]\, Y => \prdata_39_0_iv_3[15]\);
    
    \prdata_RNO_14[2]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[2]\, C
         => \delta_f2_f0_m_i[2]\, Y => \prdata_39_0_iv_4[2]\);
    
    \prdata_RNO_7[17]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[17]\, 
        C => \addr_matrix_f2_m_i[17]\, Y => 
        \prdata_39_0_iv_1[17]\);
    
    \prdata_RNO_13[1]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[1]\, 
        Y => \addr_matrix_f2_m_i[1]\);
    
    \reg_sp.addr_matrix_f0_1[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[26]\);
    
    \prdata_RNO_9[10]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[10]\, Y => \addr_matrix_f0_1_m_i[10]\);
    
    \prdata_RNO_3[13]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[13]\, 
        Y => \addr_data_f1_m_i[13]\);
    
    \prdata_RNO_7[20]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[20]\, C
         => \addr_matrix_f2_m_i[20]\, Y => \prdata_39_0_iv_1[20]\);
    
    \status_full_ack_RNO[1]\ : NOR3A
      port map(A => \status_full_0[1]\, B => apbi_c_51, C => 
        N_933_0, Y => \status_full_ack_8[1]\);
    
    \reg_wp.addr_data_f1[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[9]\);
    
    \reg_wp.addr_data_f0[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[27]\);
    
    \prdata_RNO_17[0]\ : OR2B
      port map(A => \status_full_0[0]\, B => prdata_13_sqmuxa, Y
         => \status_full_m_i[0]\);
    
    \reg_wp.delta_snapshot[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[3]\);
    
    \prdata_RNO_4[19]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[19]\, Y
         => \addr_data_f1_m_i[19]\);
    
    \prdata_RNO[14]\ : OR3C
      port map(A => \prdata_39_0_iv_2[14]\, B => 
        \delta_snapshot_m_i[14]\, C => \prdata_39_0_iv_6[14]\, Y
         => \prdata_39[14]\);
    
    \reg_wp.status_full_err_RNO_0[3]\ : NOR3A
      port map(A => N_933_0, B => \status_full_err[3]\, C => 
        status_full_err_0(3), Y => N_145);
    
    \prdata_RNO_2[30]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[30]\, B => 
        \addr_matrix_f0_0_m_i[30]\, C => \prdata_39_0_iv_1[30]\, 
        Y => \prdata_39_0_iv_4[30]\);
    
    \reg_sp.addr_matrix_f1[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[1]\);
    
    \prdata_RNO_6[27]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[27]\, 
        Y => \addr_matrix_f0_0_m_i[27]\);
    
    \prdata_RNO_3[30]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[30]\, Y
         => \addr_data_f2_m_i[30]\);
    
    \prdata_RNO_6[7]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[7]\, Y
         => \delta_f2_f0_m_i[7]\);
    
    \reg_sp.addr_matrix_f0_0[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[11]\);
    
    \reg_wp.addr_data_f3[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[14]\);
    
    \prdata_RNO_1[22]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[22]\, C
         => \addr_data_f1_m_i[22]\, Y => \prdata_39_0_iv_2[22]\);
    
    \prdata_RNO[28]\ : OR3C
      port map(A => \prdata_39_0_iv_3[28]\, B => 
        \prdata_39_0_iv_2[28]\, C => \prdata_39_0_iv_4[28]\, Y
         => \prdata_39[28]\);
    
    \prdata_RNO_4[20]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[20]\, Y
         => \addr_data_f1_m_i[20]\);
    
    \status_full_ack_RNO[3]\ : NOR3A
      port map(A => \status_full_0[3]\, B => apbi_c_53, C => 
        \status_full_5_i_o2[0]\, Y => \status_full_ack_8[3]\);
    
    \reg_wp.nb_burst_available_1_sqmuxa_0_a2_1\ : NOR3A
      port map(A => apbi_c_20, B => apbi_c_21, C => apbi_c_22, Y
         => N_159);
    
    \reg_wp.addr_data_f2[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[8]\);
    
    \prdata_RNO_14[8]\ : OR2B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[8]\, Y
         => \addr_matrix_f1_m_i[8]\);
    
    \prdata_RNO_13[7]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[7]\, 
        Y => \addr_matrix_f0_1_m_i[7]\);
    
    \reg_wp.delta_f2_f1[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[5]\);
    
    \reg_wp.nb_snapshot_param[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[5]\);
    
    \reg_wp.addr_data_f2[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[19]\);
    
    \prdata_RNO_1[18]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[18]\, C => \addr_matrix_f0_1_m_i[18]\, 
        Y => \prdata_39_0_iv_0[18]\);
    
    \reg_wp.addr_data_f0[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[17]\);
    
    \prdata_RNO_14[4]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[4]\, 
        C => \addr_matrix_f2_m_i[4]\, Y => \prdata_39_0_iv_1[4]\);
    
    \prdata_RNO_5[15]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[15]\, 
        C => \addr_matrix_f2_m_i[15]\, Y => 
        \prdata_39_0_iv_1[15]\);
    
    \reg_wp.status_full_err_RNO_0[2]\ : NOR3A
      port map(A => N_933_0, B => \status_full_err[2]\, C => 
        status_full_err_0(2), Y => N_143);
    
    \prdata_RNO_6[2]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[2]\, C
         => enable_f2_m_i, Y => \prdata_39_0_iv_7[2]\);
    
    \prdata_RNO_2[15]\ : NOR3C
      port map(A => \addr_data_f1_m_i[15]\, B => 
        \addr_data_f0_m_i[15]\, C => \delta_snapshot_m_i[15]\, Y
         => \prdata_39_0_iv_5[15]\);
    
    \prdata_RNO_8[13]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[13]\, Y => \addr_matrix_f0_1_m_i[13]\);
    
    \reg_wp.addr_data_f3[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[18]\);
    
    prdata_5_sqmuxa_0_a2_0 : NOR2A
      port map(A => N_172, B => N_157, Y => prdata_5_sqmuxa_0);
    
    \prdata_RNO_4[2]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[2]\, C
         => status_ready_matrix_f1_m_i, Y => 
        \prdata_39_0_iv_2[2]\);
    
    \prdata_RNO_2[29]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[29]\, B => 
        \addr_matrix_f0_0_m_i[29]\, C => \prdata_39_0_iv_1[29]\, 
        Y => \prdata_39_0_iv_4[29]\);
    
    \prdata_RNO_0[20]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[20]\, 
        C => \addr_data_f2_m_i[20]\, Y => \prdata_39_0_iv_3[20]\);
    
    \reg_sp.addr_matrix_f2[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[16]\);
    
    \reg_wp.delta_f2_f1[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[0]\);
    
    \prdata_RNO_15[0]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[0]\, 
        Y => \addr_data_f2_m_i[0]\);
    
    \reg_wp.status_new_err_RNO[1]\ : OA1B
      port map(A => apbi_c_59, B => \status_full_5_i_o2[0]\, C
         => N_149, Y => \status_new_err_RNO[1]\);
    
    \prdata_RNO_1[6]\ : AOI1B
      port map(A => \nb_snapshot_param[6]\, B => prdata_18_sqmuxa, 
        C => \prdata_39_0_iv_5[6]\, Y => \prdata_39_0_iv_9[6]\);
    
    \reg_sp.addr_matrix_f2[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[11]\);
    
    \reg_sp.addr_matrix_f2[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[10]\);
    
    \reg_sp.addr_matrix_f0_0[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[18]\);
    
    \prdata_RNO_20[3]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \enable_f3\, Y => 
        enable_f3_m_i);
    
    \reg_sp.addr_matrix_f0_0[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[29]\);
    
    \prdata_RNO_10[8]\ : AOI1B
      port map(A => \status_new_err[0]\, B => prdata_13_sqmuxa, C
         => \addr_data_f0_m_i[8]\, Y => \prdata_39_0_iv_2[8]\);
    
    \prdata_RNO_3[7]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[7]\, Y
         => \delta_snapshot_m_i[7]\);
    
    \reg_wp.delta_f2_f1[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[4]\);
    
    \reg_sp.addr_matrix_f0_1[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[20]\);
    
    \prdata_RNO_4[30]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[30]\, Y
         => \addr_data_f1_m_i[30]\);
    
    \reg_sp.addr_matrix_f2[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[26]\);
    
    \reg_sp.addr_matrix_f0_1[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[23]\);
    
    \prdata_RNO_5[18]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[18]\, Y
         => \addr_data_f3_m_i[18]\);
    
    \reg_wp.delta_snapshot[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[15]\);
    
    \prdata_RNO_2[18]\ : NOR3C
      port map(A => \addr_data_f3_m_i[18]\, B => 
        \addr_data_f2_m_i[18]\, C => \prdata_39_0_iv_2[18]\, Y
         => \prdata_39_0_iv_5[18]\);
    
    \reg_wp.data_shaping_R1\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => data_shaping_BW_1_sqmuxa, Q => data_shaping_R1);
    
    \prdata_RNO_12[6]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[6]\, 
        Y => \addr_matrix_f0_0_m_i[6]\);
    
    \reg_sp.addr_matrix_f0_1[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[12]\);
    
    \reg_wp.delta_snapshot[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[0]\);
    
    \reg_sp.addr_matrix_f2[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[21]\);
    
    \reg_sp.addr_matrix_f0_0_1_sqmuxa_0_a2\ : NOR3C
      port map(A => N_159, B => N_928, C => N_930, Y => 
        addr_matrix_f0_0_1_sqmuxa);
    
    \prdata_RNO_0[0]\ : NOR3C
      port map(A => \delta_snapshot_m_i[0]\, B => 
        \prdata_39_0_iv_2[0]\, C => \prdata_39_0_iv_9[0]\, Y => 
        \prdata_39_0_iv_13[0]\);
    
    \prdata_RNO_8[1]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[1]\, B => 
        \addr_matrix_f0_0_m_i[1]\, C => \status_full_m_i[1]\, Y
         => \prdata_39_0_iv_6[1]\);
    
    \reg_wp.enable_f3\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \enable_f3\);
    
    \prdata[24]\ : DFN1C0
      port map(D => \prdata_39[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(24));
    
    \prdata_RNO[22]\ : OR3C
      port map(A => \prdata_39_0_iv_3[22]\, B => 
        \prdata_39_0_iv_2[22]\, C => \prdata_39_0_iv_4[22]\, Y
         => \prdata_39[22]\);
    
    \reg_sp.addr_matrix_f2[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[20]\);
    
    \prdata_RNO_4[15]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[15]\, 
        Y => \addr_matrix_f0_0_m_i[15]\);
    
    \prdata_RNO_18[0]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[0]\, Y
         => \delta_f2_f1_m_i[0]\);
    
    \prdata_RNO_13[2]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[2]\, Y
         => \delta_f2_f1_m_i[2]\);
    
    \prdata_RNO_8[8]\ : OR2B
      port map(A => \nb_snapshot_param[8]\, B => prdata_18_sqmuxa, 
        Y => \nb_snapshot_param_m_i[8]\);
    
    \prdata_RNO_8[21]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[21]\, Y
         => \addr_data_f1_m_i[21]\);
    
    \prdata_RNO_8[26]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[26]\, Y
         => \addr_matrix_f2_m_i[26]\);
    
    \prdata_RNO_1[17]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[17]\, C
         => \addr_data_f1_m_i[17]\, Y => \prdata_39_0_iv_2[17]\);
    
    \prdata_RNO_14[9]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[9]\, 
        Y => \addr_matrix_f0_0_m_i[9]\);
    
    \prdata_RNO[20]\ : OR3C
      port map(A => \prdata_39_0_iv_3[20]\, B => 
        \prdata_39_0_iv_2[20]\, C => \prdata_39_0_iv_4[20]\, Y
         => \prdata_39[20]\);
    
    \prdata_RNO_15[5]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[5]\, Y
         => \delta_f2_f1_m_i[5]\);
    
    \prdata_RNO_12[3]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[3]\, Y
         => \addr_data_f3_m_i[3]\);
    
    \reg_sp.addr_matrix_f0_1[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[31]\);
    
    \prdata_RNO_5[24]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[24]\, 
        Y => \addr_matrix_f0_1_m_i[24]\);
    
    \reg_sp.addr_matrix_f1[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[5]\);
    
    prdata_15_sqmuxa_0_a2 : NOR2B
      port map(A => N_164, B => N_161, Y => prdata_15_sqmuxa);
    
    \reg_wp.delta_snapshot[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[12]\);
    
    \prdata_RNO_19[1]\ : AOI1B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[1]\, C
         => \delta_f2_f1_m_i[1]\, Y => \prdata_39_0_iv_5[1]\);
    
    \reg_wp.status_new_err_RNO_0[2]\ : NOR3A
      port map(A => N_933_0, B => \status_new_err[2]\, C => 
        status_new_err_0_2, Y => N_151);
    
    \prdata_RNO_6[11]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[11]\, Y
         => \addr_data_f3_m_i[11]\);
    
    \prdata_RNO_6[16]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[16]\, 
        Y => \addr_matrix_f0_0_m_i[16]\);
    
    \prdata_RNO_3[10]\ : AOI1B
      port map(A => prdata_2_sqmuxa_0, B => 
        \addr_matrix_f0_0[10]\, C => \addr_matrix_f0_1_m_i[10]\, 
        Y => \prdata_39_0_iv_0[10]\);
    
    \prdata_RNO_14[5]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[5]\, 
        C => \addr_matrix_f2_m_i[5]\, Y => \prdata_39_0_iv_1[5]\);
    
    \prdata_RNO_17[3]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[3]\, Y
         => \delta_snapshot_m_i[3]\);
    
    \prdata_RNO_8[22]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[22]\, Y
         => \addr_matrix_f2_m_i[22]\);
    
    prdata_17_sqmuxa_0_a2 : NOR3B
      port map(A => N_158, B => N_159, C => apbi_c_19, Y => 
        prdata_17_sqmuxa);
    
    \reg_sp.addr_matrix_f0_1_1_sqmuxa_0_a2_0_0\ : NOR3C
      port map(A => N_159, B => N_928, C => N_166, Y => 
        addr_matrix_f0_1_1_sqmuxa_0);
    
    \reg_wp.addr_data_f1[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[30]\);
    
    \prdata_RNO_2[25]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[25]\, B => 
        \addr_matrix_f0_0_m_i[25]\, C => \prdata_39_0_iv_1[25]\, 
        Y => \prdata_39_0_iv_4[25]\);
    
    \prdata_RNO_4[18]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[18]\, 
        Y => \addr_matrix_f0_1_m_i[18]\);
    
    \reg_wp.nb_burst_available[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[2]\);
    
    \prdata_RNO_8[6]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[6]\, 
        Y => \addr_matrix_f2_m_i[6]\);
    
    \prdata_RNO_3[3]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[3]\, C
         => \addr_data_f2_m_i[3]\, Y => \prdata_39_0_iv_3[3]\);
    
    \reg_wp.delta_snapshot[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[14]\);
    
    \reg_wp.delta_f2_f1[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f1_1_sqmuxa, Q => \delta_f2_f1[9]\);
    
    \reg_sp.addr_matrix_f2[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[14]\);
    
    \prdata_RNO_6[12]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[12]\, 
        C => \addr_data_f2_m_i[12]\, Y => \prdata_39_0_iv_3[12]\);
    
    \prdata_RNO_9[5]\ : OR2B
      port map(A => \nb_burst_available[5]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[5]\);
    
    \prdata_RNO_5[0]\ : AOI1B
      port map(A => \nb_burst_available[0]\, B => 
        prdata_17_sqmuxa, C => enable_f0_m_i, Y => 
        \prdata_39_0_iv_9[0]\);
    
    \reg_wp.addr_data_f3[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[27]\);
    
    \prdata_RNO_5[17]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[17]\, 
        Y => \addr_matrix_f0_1_m_i[17]\);
    
    \prdata_RNO_17[7]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[7]\, Y
         => \addr_data_f0_m_i[7]\);
    
    \prdata_RNO_2[17]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[17]\, B => 
        \addr_matrix_f0_0_m_i[17]\, C => \prdata_39_0_iv_1[17]\, 
        Y => \prdata_39_0_iv_4[17]\);
    
    \reg_wp.nb_snapshot_param[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[10]\);
    
    \reg_sp.addr_matrix_f1[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[16]\);
    
    \reg_wp.delta_snapshot[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[11]\);
    
    \reg_sp.config_active_interruption_onNewMatrix\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => config_active_interruption_onError_0_sqmuxa, Q => 
        config_active_interruption_onNewMatrix);
    
    \reg_wp.addr_data_f1[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[31]\);
    
    \reg_wp.status_full_RNO[3]\ : OA1B
      port map(A => apbi_c_53, B => \status_full_5_i_o2[0]\, C
         => N_138, Y => \status_full_RNO[3]\);
    
    \prdata_RNO_3[24]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[24]\, Y
         => \addr_data_f2_m_i[24]\);
    
    \reg_wp.addr_data_f3[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[19]\);
    
    \prdata_RNO_2[8]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[8]\, B => 
        \prdata_39_0_iv_2[8]\, C => \nb_burst_available_m_i[8]\, 
        Y => \prdata_39_0_iv_10[8]\);
    
    \reg_sp.addr_matrix_f1[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[11]\);
    
    \status_full_ack_RNO[2]\ : NOR3A
      port map(A => \status_full_0[2]\, B => apbi_c_52, C => 
        N_933_0, Y => \status_full_ack_8[2]\);
    
    \reg_sp.addr_matrix_f0_1[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[24]\);
    
    \reg_sp.addr_matrix_f0_1[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[3]\);
    
    \reg_sp.addr_matrix_f0_1[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => 
        \addr_matrix_f0_1[25]\);
    
    \prdata_RNO_8[10]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[10]\, 
        C => \prdata_39_0_iv_1[10]\, Y => \prdata_39_0_iv_5[10]\);
    
    \reg_sp.addr_matrix_f1[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[10]\);
    
    \reg_sp.status_error_anticipating_empty_fifo_1_sqmuxa_0_a2\ : 
        NOR3
      port map(A => N_157, B => un1_apbi_2, C => N_169, Y => 
        status_error_anticipating_empty_fifo_1_sqmuxa);
    
    prdata_3_sqmuxa_0_a2 : NOR3C
      port map(A => N_159, B => N_928, C => apbi_c_19, Y => 
        prdata_3_sqmuxa);
    
    \prdata_RNO_3[0]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[0]\, Y
         => \delta_snapshot_m_i[0]\);
    
    \prdata_RNO_2[2]\ : NOR3C
      port map(A => \prdata_39_0_iv_6[2]\, B => 
        \nb_snapshot_param_m_i[2]\, C => data_shaping_SP1_m_i, Y
         => \prdata_39_0_iv_13[2]\);
    
    \prdata_RNO_7[7]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[7]\, Y
         => \addr_data_f3_m_i[7]\);
    
    \prdata_RNO_13[5]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[5]\, 
        Y => \addr_matrix_f0_0_m_i[5]\);
    
    \prdata_RNO_3[4]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[4]\, C
         => \addr_data_f1_m_i[4]\, Y => \prdata_39_0_iv_3[4]\);
    
    \lpp_top_apbreg.un1_apbi_2\ : OR2B
      port map(A => apbi_c_49, B => apbi_c_16, Y => un1_apbi_2);
    
    \reg_wp.status_full_err_RNO[3]\ : OA1B
      port map(A => apbi_c_57, B => \status_full_5_i_o2[0]\, C
         => N_145, Y => \status_full_err_RNO[3]\);
    
    \reg_sp.addr_matrix_f2[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[7]\);
    
    \reg_sp.addr_matrix_f2[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[24]\);
    
    \reg_wp.addr_data_f1[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[24]\);
    
    \prdata_RNO_5[6]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[6]\, C
         => \addr_data_f2_m_i[6]\, Y => \prdata_39_0_iv_3[6]\);
    
    \prdata_RNO_2[28]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[28]\, B => 
        \addr_matrix_f0_0_m_i[28]\, C => \prdata_39_0_iv_1[28]\, 
        Y => \prdata_39_0_iv_4[28]\);
    
    \prdata_RNO_16[4]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => \addr_data_f2[4]\, 
        Y => \addr_data_f2_m_i[4]\);
    
    \prdata_RNO[17]\ : OR3C
      port map(A => \prdata_39_0_iv_3[17]\, B => 
        \prdata_39_0_iv_2[17]\, C => \prdata_39_0_iv_4[17]\, Y
         => \prdata_39[17]\);
    
    \reg_wp.addr_data_f0[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[23]\);
    
    \prdata_RNO[25]\ : OR3C
      port map(A => \prdata_39_0_iv_3[25]\, B => 
        \prdata_39_0_iv_2[25]\, C => \prdata_39_0_iv_4[25]\, Y
         => \prdata_39[25]\);
    
    \prdata[20]\ : DFN1C0
      port map(D => \prdata_39[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(20));
    
    \reg_wp.addr_data_f0[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[20]\);
    
    \prdata_RNO_1[4]\ : AOI1B
      port map(A => \nb_snapshot_param[4]\, B => prdata_18_sqmuxa, 
        C => \prdata_39_0_iv_6[4]\, Y => \prdata_39_0_iv_10[4]\);
    
    \prdata_RNO_21[1]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[1]\, Y
         => \delta_f2_f1_m_i[1]\);
    
    \reg_wp.addr_data_f3[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[1]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \prdata_RNO_8[3]\ : NOR3C
      port map(A => \delta_snapshot_m_i[3]\, B => 
        \prdata_39_0_iv_1[3]\, C => \nb_burst_available_m_i[3]\, 
        Y => \prdata_39_0_iv_11[3]\);
    
    \reg_sp.addr_matrix_f0_0[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[27]\);
    
    \prdata_RNO_1[29]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[29]\, C
         => \addr_data_f1_m_i[29]\, Y => \prdata_39_0_iv_2[29]\);
    
    \prdata_RNO_5[23]\ : OR2B
      port map(A => prdata_12_sqmuxa, B => \addr_data_f3[23]\, Y
         => \addr_data_f3_m_i[23]\);
    
    \prdata_RNO_17[8]\ : OR2B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[8]\, Y
         => \addr_data_f0_m_i[8]\);
    
    \prdata_RNO_10[6]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[6]\, Y
         => \delta_snapshot_m_i[6]\);
    
    \prdata_RNO_0[14]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[14]\, C
         => \addr_data_f1_m_i[14]\, Y => \prdata_39_0_iv_2[14]\);
    
    prdata_14_sqmuxa_0_a2 : NOR3B
      port map(A => apbi_c_21, B => apbi_c_19, C => N_931, Y => 
        prdata_14_sqmuxa);
    
    \reg_wp.addr_data_f1[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[28]\);
    
    \reg_wp.delta_snapshot[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[13]\);
    
    \prdata_RNO_8[7]\ : OR2B
      port map(A => \nb_snapshot_param[7]\, B => prdata_18_sqmuxa, 
        Y => \nb_snapshot_param_m_i[7]\);
    
    \reg_wp.addr_data_f0[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[21]\);
    
    prdata_3_sqmuxa_0_a2_0 : NOR3C
      port map(A => N_159, B => N_928, C => apbi_c_19, Y => 
        prdata_3_sqmuxa_0);
    
    \prdata[23]\ : DFN1C0
      port map(D => \prdata_39[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(23));
    
    \prdata_RNO_4[17]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[17]\, 
        Y => \addr_data_f1_m_i[17]\);
    
    \reg_wp.delta_f2_f0[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[6]\);
    
    \prdata_RNO_9[11]\ : AOI1B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[11]\, 
        C => \addr_data_f2_m_i[11]\, Y => \prdata_39_0_iv_3[11]\);
    
    \prdata_RNO_7[21]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[21]\, C
         => \addr_data_f1_m_i[21]\, Y => \prdata_39_0_iv_2[21]\);
    
    \prdata_RNO_7[26]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[26]\, C
         => \addr_matrix_f2_m_i[26]\, Y => \prdata_39_0_iv_1[26]\);
    
    \prdata_RNO[9]\ : OR3C
      port map(A => \prdata_39_0_iv_9[9]\, B => 
        \prdata_39_0_iv_8[9]\, C => \prdata_39_0_iv_10[9]\, Y => 
        \prdata_39[9]\);
    
    \reg_wp.addr_data_f0[13]\ : DFN1E1C0
      port map(D => apbi_c_63, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[13]\);
    
    \prdata_RNO_20[2]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[2]\, 
        Y => \addr_matrix_f2_m_i[2]\);
    
    \prdata_RNO_12[7]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[7]\, 
        Y => \addr_matrix_f2_m_i[7]\);
    
    \reg_wp.addr_data_f0[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[10]\);
    
    \prdata_RNO_2[31]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[31]\, B => 
        \addr_matrix_f0_0_m_i[31]\, C => \prdata_39_0_iv_1[31]\, 
        Y => \prdata_39_0_iv_4[31]\);
    
    \prdata_RNO_13[3]\ : AOI1B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[3]\, C
         => enable_f3_m_i, Y => \prdata_39_0_iv_5[3]\);
    
    \prdata_RNO_14[3]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => \addr_matrix_f0_1[3]\, 
        Y => \addr_matrix_f0_1_m_i[3]\);
    
    \prdata_RNO_3[31]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[31]\, Y
         => \addr_data_f2_m_i[31]\);
    
    \reg_wp.addr_data_f2_1_sqmuxa_0_a2_0\ : NOR3C
      port map(A => apbi_c_22, B => N_928, C => apbi_c_21, Y => 
        N_168);
    
    \prdata_RNO_5[5]\ : AOI1B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[5]\, C
         => \prdata_39_0_iv_2[5]\, Y => \prdata_39_0_iv_7[5]\);
    
    \reg_wp.addr_data_f1[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[14]\);
    
    \reg_sp.addr_matrix_f2[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa_0, Q => \addr_matrix_f2[1]\);
    
    \reg_wp.delta_snapshot[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_snapshot_1_sqmuxa, Q => \delta_snapshot[9]\);
    
    \prdata[30]\ : DFN1C0
      port map(D => \prdata_39[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(30));
    
    \prdata_RNO_13[8]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[8]\, 
        Y => \addr_matrix_f2_m_i[8]\);
    
    \reg_wp.status_new_err[3]\ : DFN1C0
      port map(D => \status_new_err_RNO[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_new_err_0[3]\);
    
    \reg_wp.addr_data_f1[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[0]\);
    
    \prdata_RNO_12[2]\ : OR2B
      port map(A => \status_full_0[2]\, B => prdata_13_sqmuxa, Y
         => \status_full_m_i[2]\);
    
    \reg_wp.delta_f2_f0[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => delta_f2_f0_1_sqmuxa, Q => \delta_f2_f0[4]\);
    
    \prdata_RNO_12[1]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \enable_f1\, Y => 
        enable_f1_m_i);
    
    \prdata[11]\ : DFN1C0
      port map(D => \prdata_39[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(11));
    
    \reg_sp.addr_matrix_f0_0[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[19]\);
    
    \reg_wp.addr_data_f2_1_sqmuxa_0_a2_0_0\ : NOR3C
      port map(A => apbi_c_22, B => N_928, C => apbi_c_21, Y => 
        N_168_0);
    
    \reg_wp.addr_data_f0[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[11]\);
    
    \prdata_RNO_4[21]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[21]\, 
        Y => \addr_matrix_f0_1_m_i[21]\);
    
    \prdata_RNO_4[26]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[26]\, Y
         => \addr_data_f1_m_i[26]\);
    
    \prdata_RNO_9[12]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[12]\, Y => \addr_data_f2_m_i[12]\);
    
    \prdata_RNO_3[23]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[23]\, Y
         => \addr_matrix_f2_m_i[23]\);
    
    \prdata_RNO_7[22]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[22]\, C
         => \addr_matrix_f2_m_i[22]\, Y => \prdata_39_0_iv_1[22]\);
    
    \reg_sp.addr_matrix_f0_1[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[5]\);
    
    \reg_wp.addr_data_f1[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[18]\);
    
    \prdata_RNO_2[27]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[27]\, B => 
        \addr_matrix_f0_0_m_i[27]\, C => \prdata_39_0_iv_1[27]\, 
        Y => \prdata_39_0_iv_4[27]\);
    
    \prdata_RNO_9[0]\ : NOR3C
      port map(A => \status_full_m_i[0]\, B => 
        \delta_f2_f1_m_i[0]\, C => \prdata_39_0_iv_5[0]\, Y => 
        \prdata_39_0_iv_11[0]\);
    
    \reg_sp.status_ready_matrix_f0_1\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_ready_matrix_f0_1);
    
    \reg_sp.addr_matrix_f1[14]\ : DFN1E1C0
      port map(D => apbi_c_64, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[14]\);
    
    \prdata_RNO_5[8]\ : NOR3C
      port map(A => \addr_matrix_f2_m_i[8]\, B => 
        \addr_matrix_f1_m_i[8]\, C => \delta_snapshot_m_i[8]\, Y
         => \prdata_39_0_iv_6[8]\);
    
    \prdata_RNO[30]\ : OR3C
      port map(A => \prdata_39_0_iv_3[30]\, B => 
        \prdata_39_0_iv_2[30]\, C => \prdata_39_0_iv_4[30]\, Y
         => \prdata_39[30]\);
    
    \apbo.pirq_RNO_2[15]\ : NOR3A
      port map(A => \pirq_2_i_a2_5[15]\, B => status_full(1), C
         => status_full(0), Y => \pirq_2_i_a2_8[15]\);
    
    \prdata_RNO_0[21]\ : AOI1B
      port map(A => prdata_4_sqmuxa, B => \addr_matrix_f1[21]\, C
         => \addr_matrix_f2_m_i[21]\, Y => \prdata_39_0_iv_1[21]\);
    
    \reg_sp.addr_matrix_f0_1[11]\ : DFN1E1C0
      port map(D => apbi_c_61, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[11]\);
    
    \prdata_RNO_7[14]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[14]\, 
        Y => \addr_matrix_f2_m_i[14]\);
    
    \prdata_RNO_11[0]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \enable_f0\, Y => 
        enable_f0_m_i);
    
    \prdata_RNO_0[26]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[26]\, 
        C => \addr_data_f2_m_i[26]\, Y => \prdata_39_0_iv_3[26]\);
    
    \prdata_RNO_4[8]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[8]\, Y
         => \delta_f2_f1_m_i[8]\);
    
    \reg_sp.addr_matrix_f0_0[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[5]\);
    
    prdata_12_sqmuxa_0_a2 : NOR2A
      port map(A => N_168, B => N_157, Y => prdata_12_sqmuxa);
    
    \prdata_RNO_21[3]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[3]\, 
        Y => \addr_matrix_f2_m_i[3]\);
    
    \prdata_RNO_4[22]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[22]\, Y
         => \addr_data_f1_m_i[22]\);
    
    \reg_wp.addr_data_f0[9]\ : DFN1E1C0
      port map(D => apbi_c_59, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[9]\);
    
    prdata_5_sqmuxa_0_a2 : NOR2A
      port map(A => N_172, B => N_157, Y => prdata_5_sqmuxa);
    
    \reg_wp.addr_data_f2[2]\ : DFN1E1C0
      port map(D => apbi_c_52, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[2]\);
    
    \prdata_RNO_6[30]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[30]\, 
        Y => \addr_matrix_f0_0_m_i[30]\);
    
    \prdata_RNO_6[24]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[24]\, 
        Y => \addr_matrix_f0_0_m_i[24]\);
    
    \reg_sp.addr_matrix_f1_1_sqmuxa_0_a2_1\ : NOR3B
      port map(A => apbi_c_21, B => N_928, C => apbi_c_22, Y => 
        N_172);
    
    \reg_wp.addr_data_f0[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[25]\);
    
    \reg_sp.addr_matrix_f0_0[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => \addr_matrix_f0_0[7]\);
    
    \prdata_RNO_17[2]\ : OR2B
      port map(A => prdata_2_sqmuxa_0, B => \addr_matrix_f0_0[2]\, 
        Y => \addr_matrix_f0_0_m_i[2]\);
    
    \prdata_RNO_0[13]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[13]\, C
         => \addr_data_f1_m_i[13]\, Y => \prdata_39_0_iv_2[13]\);
    
    \reg_wp.nb_snapshot_param[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[8]\);
    
    \reg_wp.addr_data_f0[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa, Q => \addr_data_f0[26]\);
    
    \reg_sp.addr_matrix_f2_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_172, B => N_157, C => un1_apbi_2, Y => 
        addr_matrix_f2_1_sqmuxa);
    
    \reg_wp.delta_snapshot_1_sqmuxa_0_a2\ : NOR3B
      port map(A => apbi_c_21, B => N_166, C => N_931, Y => 
        delta_snapshot_1_sqmuxa);
    
    \reg_sp.addr_matrix_f0_1[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa, Q => \addr_matrix_f0_1[6]\);
    
    \prdata_RNO_1[25]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[25]\, C
         => \addr_data_f1_m_i[25]\, Y => \prdata_39_0_iv_2[25]\);
    
    \reg_wp.addr_data_f1_1_sqmuxa_0_a2_0\ : NOR3A
      port map(A => N_166, B => apbi_c_21, C => N_931, Y => 
        addr_data_f1_1_sqmuxa_0);
    
    \prdata_RNO_15[1]\ : AOI1B
      port map(A => prdata_0_sqmuxa, B => 
        config_active_interruption_onError, C => 
        status_ready_matrix_f0_1_m_i, Y => \prdata_39_0_iv_2[1]\);
    
    \reg_wp.addr_data_f2[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa_0, Q => \addr_data_f2[17]\);
    
    \prdata_RNO[11]\ : OR3C
      port map(A => \prdata_39_0_iv_5[11]\, B => 
        \prdata_39_0_iv_4[11]\, C => \prdata_39_0_iv_6[11]\, Y
         => \prdata_39[11]\);
    
    \prdata[25]\ : DFN1C0
      port map(D => \prdata_39[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(25));
    
    \prdata_RNO_1[8]\ : NOR3C
      port map(A => \delta_f2_f0_m_i[8]\, B => 
        \addr_data_f3_m_i[8]\, C => \nb_snapshot_param_m_i[8]\, Y
         => \prdata_39_0_iv_8[8]\);
    
    \prdata_RNO_0[22]\ : AOI1B
      port map(A => prdata_12_sqmuxa_0, B => \addr_data_f3[22]\, 
        C => \addr_data_f2_m_i[22]\, Y => \prdata_39_0_iv_3[22]\);
    
    \prdata_RNO_4[31]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[31]\, Y
         => \addr_data_f1_m_i[31]\);
    
    \reg_wp.addr_data_f2[24]\ : DFN1E1C0
      port map(D => apbi_c_74, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[24]\);
    
    \reg_wp.status_full_err_RNO_0[1]\ : NOR3A
      port map(A => N_933_0, B => \status_full_err[1]\, C => 
        status_full_err_0(1), Y => N_141);
    
    \reg_sp.addr_matrix_f2_1_sqmuxa_0_a2_0\ : NOR3A
      port map(A => N_172, B => N_157, C => un1_apbi_2, Y => 
        addr_matrix_f2_1_sqmuxa_0);
    
    \reg_sp.addr_matrix_f2[8]\ : DFN1E1C0
      port map(D => apbi_c_58, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[8]\);
    
    \prdata_RNO_8[9]\ : OR2B
      port map(A => \nb_snapshot_param[9]\, B => prdata_18_sqmuxa, 
        Y => \nb_snapshot_param_m_i[9]\);
    
    \status_full_ack[3]\ : DFN1C0
      port map(D => \status_full_ack_8[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => status_full_ack(3));
    
    \reg_wp.delta_f2_f0_1_sqmuxa_0_a2\ : NOR3A
      port map(A => N_164, B => N_157, C => un1_apbi_2, Y => 
        delta_f2_f0_1_sqmuxa);
    
    \prdata_RNO[29]\ : OR3C
      port map(A => \prdata_39_0_iv_3[29]\, B => 
        \prdata_39_0_iv_2[29]\, C => \prdata_39_0_iv_4[29]\, Y
         => \prdata_39[29]\);
    
    \prdata_RNO_14[0]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[0]\, 
        C => \addr_matrix_f2_m_i[0]\, Y => \prdata_39_0_iv_1[0]\);
    
    \prdata_RNO_6[5]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[5]\, B => 
        \addr_matrix_f0_0_m_i[5]\, C => \prdata_39_0_iv_1[5]\, Y
         => \prdata_39_0_iv_6[5]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \prdata_RNO_8[29]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[29]\, Y
         => \addr_matrix_f2_m_i[29]\);
    
    \reg_wp.status_full[0]\ : DFN1C0
      port map(D => \status_full_RNO[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \status_full_0[0]\);
    
    \reg_sp.addr_matrix_f0_1[18]\ : DFN1E1C0
      port map(D => apbi_c_68, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_1_1_sqmuxa_0, Q => 
        \addr_matrix_f0_1[18]\);
    
    \prdata_RNO[16]\ : OR3C
      port map(A => \prdata_39_0_iv_3[16]\, B => 
        \prdata_39_0_iv_2[16]\, C => \prdata_39_0_iv_4[16]\, Y
         => \prdata_39[16]\);
    
    \prdata[0]\ : DFN1C0
      port map(D => \prdata_39[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(0));
    
    \apbo.pirq_RNO_5[15]\ : NOR2
      port map(A => status_full(2), B => status_full(3), Y => 
        \pirq_2_i_a2_5[15]\);
    
    \reg_wp.addr_data_f0_1_sqmuxa_0_a2_0\ : NOR3A
      port map(A => N_930, B => apbi_c_21, C => N_931, Y => 
        addr_data_f0_1_sqmuxa_0);
    
    \reg_wp.addr_data_f0[15]\ : DFN1E1C0
      port map(D => apbi_c_65, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[15]\);
    
    prdata_9_sqmuxa_0_a2_0 : NOR3
      port map(A => apbi_c_21, B => N_931, C => apbi_c_19, Y => 
        prdata_9_sqmuxa_0);
    
    \reg_wp.addr_data_f3[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[6]\);
    
    \reg_wp.addr_data_f2[28]\ : DFN1E1C0
      port map(D => apbi_c_78, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[28]\);
    
    \reg_wp.addr_data_f0[16]\ : DFN1E1C0
      port map(D => apbi_c_66, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[16]\);
    
    \reg_wp.status_full_err[1]\ : DFN1C0
      port map(D => \status_full_err_RNO[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \status_full_err[1]\);
    
    \reg_wp.nb_burst_available[10]\ : DFN1E1C0
      port map(D => apbi_c_60, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[10]\);
    
    \reg_wp.nb_snapshot_param[1]\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[1]\);
    
    \reg_wp.addr_data_f1[29]\ : DFN1E1C0
      port map(D => apbi_c_79, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[29]\);
    
    \reg_sp.addr_matrix_f0_0[26]\ : DFN1E1C0
      port map(D => apbi_c_76, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa, Q => 
        \addr_matrix_f0_0[26]\);
    
    \prdata_RNO_7[4]\ : OR2B
      port map(A => \nb_burst_available[4]\, B => 
        prdata_17_sqmuxa, Y => \nb_burst_available_m_i[4]\);
    
    \prdata_RNO_5[20]\ : OR2B
      port map(A => prdata_3_sqmuxa, B => \addr_matrix_f0_1[20]\, 
        Y => \addr_matrix_f0_1_m_i[20]\);
    
    \prdata_RNO_6[19]\ : OR2B
      port map(A => prdata_2_sqmuxa, B => \addr_matrix_f0_0[19]\, 
        Y => \addr_matrix_f0_0_m_i[19]\);
    
    prdata_1_sqmuxa_0_a2_0 : OR2A
      port map(A => apbi_c_19, B => apbi_c_20, Y => N_157);
    
    \reg_wp.delta_f2_f1_1_sqmuxa_0_a2\ : NOR3B
      port map(A => N_930, B => N_164, C => apbi_c_20, Y => 
        delta_f2_f1_1_sqmuxa);
    
    \reg_wp.addr_data_f2[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f2_1_sqmuxa, Q => \addr_data_f2[5]\);
    
    \reg_sp.addr_matrix_f1[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[3]\);
    
    \prdata_RNO_1[28]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[28]\, C
         => \addr_data_f1_m_i[28]\, Y => \prdata_39_0_iv_2[28]\);
    
    \reg_sp.addr_matrix_f1[25]\ : DFN1E1C0
      port map(D => apbi_c_75, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[25]\);
    
    \prdata_RNO_16[0]\ : OR2B
      port map(A => prdata_10_sqmuxa, B => \addr_data_f1[0]\, Y
         => \addr_data_f1_m_i[0]\);
    
    \reg_wp.addr_data_f3[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[23]\);
    
    \reg_wp.addr_data_f3[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[20]\);
    
    \reg_wp.nb_burst_available[0]\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[0]\);
    
    \prdata_RNO_3[11]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[11]\, 
        C => \addr_matrix_f2_m_i[11]\, Y => 
        \prdata_39_0_iv_1[11]\);
    
    \prdata_RNO_3[16]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[16]\, Y => \addr_data_f2_m_i[16]\);
    
    \reg_wp.addr_data_f3[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa, Q => \addr_data_f3[4]\);
    
    \reg_sp.addr_matrix_f1[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa_0, Q => \addr_matrix_f1[22]\);
    
    \prdata_RNO_4[4]\ : OR2B
      port map(A => prdata_8_sqmuxa, B => \burst_f0\, Y => 
        burst_f0_m_i);
    
    \prdata_RNO_7[13]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[13]\, 
        Y => \addr_matrix_f2_m_i[13]\);
    
    \prdata[9]\ : DFN1C0
      port map(D => \prdata_39[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(9));
    
    \prdata[8]\ : DFN1C0
      port map(D => \prdata_39[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(8));
    
    \prdata_RNO_10[3]\ : OR3A
      port map(A => status_ready_matrix_f2, B => N_157, C => 
        N_169, Y => status_ready_matrix_f2_m_i);
    
    \reg_sp.addr_matrix_f1[27]\ : DFN1E1C0
      port map(D => apbi_c_77, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[27]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \reg_wp.addr_data_f3[21]\ : DFN1E1C0
      port map(D => apbi_c_71, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f3_1_sqmuxa_0, Q => \addr_data_f3[21]\);
    
    \prdata_RNO_6[23]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[23]\, Y
         => \addr_data_f2_m_i[23]\);
    
    \prdata_RNO_18[5]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[5]\, 
        Y => \addr_matrix_f2_m_i[5]\);
    
    \reg_wp.addr_data_f0[22]\ : DFN1E1C0
      port map(D => apbi_c_72, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[22]\);
    
    \prdata[22]\ : DFN1C0
      port map(D => \prdata_39[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(22));
    
    \prdata_RNO_5[3]\ : NOR3C
      port map(A => \delta_f2_f0_m_i[3]\, B => 
        \addr_data_f3_m_i[3]\, C => \prdata_39_0_iv_5[3]\, Y => 
        \prdata_39_0_iv_9[3]\);
    
    \prdata_RNO_11[5]\ : AOI1B
      port map(A => \status_full_err[1]\, B => prdata_13_sqmuxa, 
        C => status_error_bad_component_error_m_i, Y => 
        \prdata_39_0_iv_2[5]\);
    
    \reg_sp.addr_matrix_f0_0[17]\ : DFN1E1C0
      port map(D => apbi_c_67, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[17]\);
    
    prdata_10_sqmuxa_0_a2 : NOR3A
      port map(A => apbi_c_19, B => apbi_c_21, C => N_931, Y => 
        prdata_10_sqmuxa);
    
    \prdata[29]\ : DFN1C0
      port map(D => \prdata_39[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(29));
    
    \prdata_RNO_4[6]\ : NOR3C
      port map(A => \addr_matrix_f0_1_m_i[6]\, B => 
        \addr_matrix_f0_0_m_i[6]\, C => \delta_f2_f1_m_i[6]\, Y
         => \prdata_39_0_iv_5[6]\);
    
    \reg_wp.nb_snapshot_param[4]\ : DFN1E1C0
      port map(D => apbi_c_54, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[4]\);
    
    \reg_wp.nb_snapshot_param[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_snapshot_param_1_sqmuxa, Q => 
        \nb_snapshot_param[7]\);
    
    \reg_wp.addr_data_f1[19]\ : DFN1E1C0
      port map(D => apbi_c_69, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa_0, Q => \addr_data_f1[19]\);
    
    \prdata_RNO_3[20]\ : OR3C
      port map(A => N_161, B => N_168, C => \addr_data_f2[20]\, Y
         => \addr_data_f2_m_i[20]\);
    
    \prdata_RNO_3[12]\ : OR2B
      port map(A => prdata_10_sqmuxa_0, B => \addr_data_f1[12]\, 
        Y => \addr_data_f1_m_i[12]\);
    
    \reg_sp.addr_matrix_f2[5]\ : DFN1E1C0
      port map(D => apbi_c_55, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f2_1_sqmuxa, Q => \addr_matrix_f2[5]\);
    
    \prdata_RNO_9[4]\ : OR3B
      port map(A => N_161_0, B => \data_shaping_R1_0\, C => N_163, 
        Y => data_shaping_R1_m_i);
    
    \prdata_RNO[4]\ : OR3C
      port map(A => \prdata_39_0_iv_11[4]\, B => 
        \prdata_39_0_iv_10[4]\, C => \prdata_39_0_iv_14[4]\, Y
         => \prdata_39[4]\);
    
    \prdata_RNO_1[14]\ : OR2B
      port map(A => prdata_14_sqmuxa, B => \delta_snapshot[14]\, 
        Y => \delta_snapshot_m_i[14]\);
    
    \prdata_RNO_6[9]\ : OR2B
      port map(A => prdata_16_sqmuxa, B => \delta_f2_f0[9]\, Y
         => \delta_f2_f0_m_i[9]\);
    
    \reg_sp.addr_matrix_f1[31]\ : DFN1E1C0
      port map(D => apbi_c_81, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[31]\);
    
    \prdata_RNO_4[1]\ : AOI1B
      port map(A => prdata_9_sqmuxa_0, B => \addr_data_f0[1]\, C
         => \addr_data_f1_m_i[1]\, Y => \prdata_39_0_iv_3[1]\);
    
    \reg_wp.nb_burst_available[3]\ : DFN1E1C0
      port map(D => apbi_c_53, CLK => HCLK_c, CLR => HRESETn_c, E
         => nb_burst_available_1_sqmuxa, Q => 
        \nb_burst_available[3]\);
    
    \reg_sp.addr_matrix_f1[30]\ : DFN1E1C0
      port map(D => apbi_c_80, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f1_1_sqmuxa, Q => \addr_matrix_f1[30]\);
    
    \prdata_RNO_8[11]\ : OR2B
      port map(A => \status_new_err_0[3]\, B => prdata_13_sqmuxa, 
        Y => \status_new_err_m_i[3]\);
    
    \prdata_RNO_8[16]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[16]\, 
        Y => \addr_matrix_f2_m_i[16]\);
    
    \reg_wp.nb_burst_available_1_sqmuxa_0_a2\ : NOR3C
      port map(A => N_158, B => N_159, C => N_930, Y => 
        nb_burst_available_1_sqmuxa);
    
    \reg_sp.status_ready_matrix_f0_0\ : DFN1E1C0
      port map(D => apbi_c_50, CLK => HCLK_c, CLR => HRESETn_c, E
         => status_error_anticipating_empty_fifo_1_sqmuxa, Q => 
        status_ready_matrix_f0_0);
    
    \prdata_RNO_0[2]\ : NOR3C
      port map(A => \prdata_39_0_iv_3[2]\, B => 
        \prdata_39_0_iv_2[2]\, C => \prdata_39_0_iv_9[2]\, Y => 
        \prdata_39_0_iv_12[2]\);
    
    \reg_wp.addr_data_f1[6]\ : DFN1E1C0
      port map(D => apbi_c_56, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[6]\);
    
    \prdata_RNO_10[10]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[10]\, Y => \addr_data_f2_m_i[10]\);
    
    \reg_wp.addr_data_f1[7]\ : DFN1E1C0
      port map(D => apbi_c_57, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f1_1_sqmuxa, Q => \addr_data_f1[7]\);
    
    \reg_wp.addr_data_f0[12]\ : DFN1E1C0
      port map(D => apbi_c_62, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_data_f0_1_sqmuxa_0, Q => \addr_data_f0[12]\);
    
    \prdata_RNO_8[25]\ : OR2B
      port map(A => prdata_5_sqmuxa, B => \addr_matrix_f2[25]\, Y
         => \addr_matrix_f2_m_i[25]\);
    
    \prdata_RNO_1[27]\ : AOI1B
      port map(A => prdata_9_sqmuxa, B => \addr_data_f0[27]\, C
         => \addr_data_f1_m_i[27]\, Y => \prdata_39_0_iv_2[27]\);
    
    \reg_sp.addr_matrix_f0_0[20]\ : DFN1E1C0
      port map(D => apbi_c_70, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[20]\);
    
    \prdata_RNO_18[4]\ : OR3A
      port map(A => status_error_anticipating_empty_fifo, B => 
        N_157, C => N_169, Y => 
        status_error_anticipating_empty_fifo_m_i);
    
    \prdata_RNO_20[4]\ : OR2B
      port map(A => prdata_15_sqmuxa, B => \delta_f2_f1[4]\, Y
         => \delta_f2_f1_m_i[4]\);
    
    \prdata_RNO_0[10]\ : NOR3C
      port map(A => \prdata_39_0_iv_0[10]\, B => 
        \addr_data_f3_m_i[10]\, C => \prdata_39_0_iv_3[10]\, Y
         => \prdata_39_0_iv_7[10]\);
    
    \reg_wp.nb_snapshot_param_1_sqmuxa_0_a2\ : NOR3C
      port map(A => N_158, B => N_159, C => N_166, Y => 
        nb_snapshot_param_1_sqmuxa);
    
    \reg_wp.enable_f1\ : DFN1E1C0
      port map(D => apbi_c_51, CLK => HCLK_c, CLR => HRESETn_c, E
         => burst_f0_1_sqmuxa, Q => \enable_f1\);
    
    \reg_sp.addr_matrix_f0_0[23]\ : DFN1E1C0
      port map(D => apbi_c_73, CLK => HCLK_c, CLR => HRESETn_c, E
         => addr_matrix_f0_0_1_sqmuxa_0, Q => 
        \addr_matrix_f0_0[23]\);
    
    \prdata_RNO_4[9]\ : AOI1B
      port map(A => prdata_4_sqmuxa_0, B => \addr_matrix_f1[9]\, 
        C => \addr_matrix_f2_m_i[9]\, Y => \prdata_39_0_iv_1[9]\);
    
    \prdata_RNO_10[15]\ : OR2B
      port map(A => prdata_5_sqmuxa_0, B => \addr_matrix_f2[15]\, 
        Y => \addr_matrix_f2_m_i[15]\);
    
    \prdata_RNO_8[12]\ : OR2B
      port map(A => prdata_3_sqmuxa_0, B => 
        \addr_matrix_f0_1[12]\, Y => \addr_matrix_f0_1_m_i[12]\);
    
    \prdata[4]\ : DFN1C0
      port map(D => \prdata_39[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => prdata_c(4));
    
    \prdata_RNO_6[15]\ : OR3C
      port map(A => N_161_0, B => N_168_0, C => 
        \addr_data_f2[15]\, Y => \addr_data_f2_m_i[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MUXN_9_2 is

    port( S_0_18          : in    std_logic;
          S_0_0           : in    std_logic;
          S_i             : in    std_logic_vector(1 to 1);
          alu_sel_coeff_0 : in    std_logic_vector(2 to 2);
          S_25            : in    std_logic;
          S_7             : in    std_logic;
          S_6             : in    std_logic;
          S_15            : in    std_logic;
          S_20            : in    std_logic;
          S_11            : in    std_logic;
          S_17            : in    std_logic;
          S_10            : in    std_logic;
          S_9             : in    std_logic;
          S_13            : in    std_logic;
          S_26            : in    std_logic;
          S_16            : in    std_logic;
          S_19            : in    std_logic;
          S_0_d0          : in    std_logic;
          S_33            : in    std_logic;
          S_12            : in    std_logic;
          S_8             : in    std_logic;
          S_22            : in    std_logic;
          S_2             : in    std_logic;
          S_23            : in    std_logic;
          S_5             : in    std_logic;
          alu_sel_coeff   : in    std_logic_vector(4 downto 3);
          alu_coef_s      : out   std_logic_vector(8 downto 0)
        );

end MUXN_9_2;

architecture DEF_ARCH of MUXN_9_2 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_43, N_19, N_47, N_25, N_48, N_28, N_49, N_50, N_56, 
        N_40, N_37, N_16, N_55, N_52, N_53, N_44, N_45, N_42, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \NB_STAGE_2.all_input.6.RES_8_1[6]\ : MX2
      port map(A => S_2, B => S_20, S => alu_sel_coeff(4), Y => 
        N_52);
    
    \NB_STAGE_2.all_input.7.RES_6_3[7]\ : MX2
      port map(A => N_55, B => N_37, S => alu_sel_coeff(3), Y => 
        alu_coef_s(7));
    
    \NB_STAGE_2.all_input.7.RES_6_2[7]\ : NOR2
      port map(A => alu_sel_coeff(4), B => S_10, Y => N_37);
    
    \NB_STAGE_2.all_input.4.RES_12_1[4]\ : MX2C
      port map(A => S_2, B => S_22, S => alu_sel_coeff(4), Y => 
        N_48);
    
    \NB_STAGE_2.all_input.0.RES_20_2[0]\ : NOR2
      port map(A => alu_sel_coeff(4), B => S_17, Y => N_16);
    
    \NB_STAGE_2.all_input.2.RES_16_2[2]\ : MX2C
      port map(A => S_15, B => S_33, S => alu_sel_coeff(4), Y => 
        N_45);
    
    \NB_STAGE_2.all_input.1.RES_18_1[1]\ : MX2C
      port map(A => S_7, B => S_25, S => alu_sel_coeff(4), Y => 
        N_43);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \NB_STAGE_2.all_input.2.RES_16_3[2]\ : MX2
      port map(A => N_44, B => N_45, S => alu_sel_coeff(3), Y => 
        alu_coef_s(2));
    
    \NB_STAGE_2.all_input.2.RES_16_1[2]\ : MX2
      port map(A => S_6, B => S_11, S => alu_sel_coeff(4), Y => 
        N_44);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \NB_STAGE_2.all_input.6.RES_8_2[6]\ : MX2C
      port map(A => S_11, B => S_33, S => alu_sel_coeff(4), Y => 
        N_53);
    
    \NB_STAGE_2.all_input.3.RES_14_1[3]\ : MX2C
      port map(A => S_5, B => S_23, S => alu_sel_coeff(4), Y => 
        N_47);
    
    \NB_STAGE_2.all_input.3.RES_14_2[3]\ : OA1C
      port map(A => S_26, B => alu_sel_coeff_0(2), C => 
        alu_sel_coeff(4), Y => N_25);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \NB_STAGE_2.all_input.3.RES_14_3[3]\ : MX2
      port map(A => N_47, B => N_25, S => alu_sel_coeff(3), Y => 
        alu_coef_s(3));
    
    \NB_STAGE_2.all_input.8.RES_4_3[8]\ : MX2
      port map(A => N_56, B => N_40, S => alu_sel_coeff(3), Y => 
        alu_coef_s(8));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \NB_STAGE_2.all_input.1.RES_18_3[1]\ : MX2
      port map(A => N_43, B => N_19, S => alu_sel_coeff(3), Y => 
        alu_coef_s(1));
    
    \NB_STAGE_2.all_input.6.RES_8_3[6]\ : MX2
      port map(A => N_52, B => N_53, S => alu_sel_coeff(3), Y => 
        alu_coef_s(6));
    
    \NB_STAGE_2.all_input.8.RES_4_1[8]\ : MX2C
      port map(A => S_0_d0, B => S_19, S => alu_sel_coeff(4), Y
         => N_56);
    
    \NB_STAGE_2.all_input.4.RES_12_3[4]\ : MX2
      port map(A => N_48, B => N_28, S => alu_sel_coeff(3), Y => 
        alu_coef_s(4));
    
    \NB_STAGE_2.all_input.4.RES_12_2[4]\ : NOR2
      port map(A => alu_sel_coeff(4), B => S_13, Y => N_28);
    
    \NB_STAGE_2.all_input.0.RES_20_3[0]\ : MX2
      port map(A => N_42, B => N_16, S => alu_sel_coeff(3), Y => 
        alu_coef_s(0));
    
    \NB_STAGE_2.all_input.8.RES_4_2[8]\ : NOR2
      port map(A => alu_sel_coeff(4), B => S_9, Y => N_40);
    
    \NB_STAGE_2.all_input.7.RES_6_1[7]\ : MX2C
      port map(A => S_i(1), B => S_19, S => alu_sel_coeff(4), Y
         => N_55);
    
    \NB_STAGE_2.all_input.1.RES_18_2[1]\ : NOR2
      port map(A => alu_sel_coeff(4), B => S_16, Y => N_19);
    
    \NB_STAGE_2.all_input.5.RES_10_1[5]\ : MX2C
      port map(A => S_5, B => S_8, S => alu_sel_coeff(4), Y => 
        N_49);
    
    \NB_STAGE_2.all_input.5.RES_10_2[5]\ : MX2C
      port map(A => S_12, B => S_33, S => alu_sel_coeff(4), Y => 
        N_50);
    
    \NB_STAGE_2.all_input.5.RES_10_3[5]\ : MX2
      port map(A => N_49, B => N_50, S => alu_sel_coeff(3), Y => 
        alu_coef_s(5));
    
    \NB_STAGE_2.all_input.0.RES_20_1[0]\ : MX2C
      port map(A => S_0_0, B => S_0_18, S => alu_sel_coeff(4), Y
         => N_42);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MUXN_9_3 is

    port( alu_coef_s        : out   std_logic_vector(8 downto 0);
          S_0_0             : in    std_logic;
          S_0_18            : in    std_logic;
          alu_sel_coeff_0_0 : in    std_logic;
          alu_sel_coeff_0_2 : in    std_logic;
          alu_sel_coeff     : in    std_logic_vector(4 downto 0)
        );

end MUXN_9_3;

architecture DEF_ARCH of MUXN_9_3 is 

  component MUXN_9_2
    port( S_0_18          : in    std_logic := 'U';
          S_0_0           : in    std_logic := 'U';
          S_i             : in    std_logic_vector(1 to 1) := (others => 'U');
          alu_sel_coeff_0 : in    std_logic_vector(2 to 2) := (others => 'U');
          S_25            : in    std_logic := 'U';
          S_7             : in    std_logic := 'U';
          S_6             : in    std_logic := 'U';
          S_15            : in    std_logic := 'U';
          S_20            : in    std_logic := 'U';
          S_11            : in    std_logic := 'U';
          S_17            : in    std_logic := 'U';
          S_10            : in    std_logic := 'U';
          S_9             : in    std_logic := 'U';
          S_13            : in    std_logic := 'U';
          S_26            : in    std_logic := 'U';
          S_16            : in    std_logic := 'U';
          S_19            : in    std_logic := 'U';
          S_0_d0          : in    std_logic := 'U';
          S_33            : in    std_logic := 'U';
          S_12            : in    std_logic := 'U';
          S_8             : in    std_logic := 'U';
          S_22            : in    std_logic := 'U';
          S_2             : in    std_logic := 'U';
          S_23            : in    std_logic := 'U';
          S_5             : in    std_logic := 'U';
          alu_sel_coeff   : in    std_logic_vector(4 downto 3) := (others => 'U');
          alu_coef_s      : out   std_logic_vector(8 downto 0)
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO14
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AXO5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI4
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AO16
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO17
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \S[0]_net_1\, \S[9]_net_1\, \S[13]_net_1\, 
        \S[16]_net_1\, \S[22]_net_1\, \S[26]_net_1\, \S[33]\, 
        \S[23]_net_1\, \S_i[1]\, \S[5]\, \S[19]\, \S[12]_net_1\, 
        \S[2]_net_1\, \S[20]_net_1\, \S[17]_net_1\, \S[10]_net_1\, 
        \S[25]_net_1\, \S[15]_net_1\, \S[11]_net_1\, \S[8]_net_1\, 
        \S[7]_net_1\, \S[6]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : MUXN_9_2
	Use entity work.MUXN_9_2(DEF_ARCH);
begin 


    \NB_STAGE_PLUS.MUXN_1\ : MUXN_9_2
      port map(S_0_18 => \S[26]_net_1\, S_0_0 => \S[8]_net_1\, 
        S_i(1) => \S_i[1]\, alu_sel_coeff_0(2) => 
        alu_sel_coeff_0_2, S_25 => \S[25]_net_1\, S_7 => 
        \S[7]_net_1\, S_6 => \S[6]_net_1\, S_15 => \S[15]_net_1\, 
        S_20 => \S[20]_net_1\, S_11 => \S[11]_net_1\, S_17 => 
        \S[17]_net_1\, S_10 => \S[10]_net_1\, S_9 => \S[9]_net_1\, 
        S_13 => \S[13]_net_1\, S_26 => S_0_18, S_16 => 
        \S[16]_net_1\, S_19 => \S[19]\, S_0_d0 => \S[0]_net_1\, 
        S_33 => \S[33]\, S_12 => \S[12]_net_1\, S_8 => S_0_0, 
        S_22 => \S[22]_net_1\, S_2 => \S[2]_net_1\, S_23 => 
        \S[23]_net_1\, S_5 => \S[5]\, alu_sel_coeff(4) => 
        alu_sel_coeff(4), alu_sel_coeff(3) => alu_sel_coeff(3), 
        alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0));
    
    \S[26]\ : AX1B
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff_0_2, C
         => alu_sel_coeff_0_0, Y => \S[26]_net_1\);
    
    \S[13]\ : XO1A
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff_0_2, C
         => alu_sel_coeff_0_0, Y => \S[13]_net_1\);
    
    \S[3]\ : XA1
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff_0_2, C
         => alu_sel_coeff(1), Y => \S[5]\);
    
    \S[9]\ : AO14
      port map(A => alu_sel_coeff_0_2, B => alu_sel_coeff(1), C
         => alu_sel_coeff_0_0, Y => \S[9]_net_1\);
    
    \S[23]\ : XA1C
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff_0_0, C
         => alu_sel_coeff_0_2, Y => \S[23]_net_1\);
    
    \S[15]\ : AXOI5
      port map(A => alu_sel_coeff(2), B => alu_sel_coeff(1), C
         => alu_sel_coeff(0), Y => \S[15]_net_1\);
    
    \S[11]\ : XAI1
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(2), C
         => alu_sel_coeff(0), Y => \S[11]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \S[8]\ : AXO5
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(0), C
         => alu_sel_coeff(2), Y => \S[8]_net_1\);
    
    \S[6]\ : AXOI4
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(0), C
         => alu_sel_coeff(2), Y => \S[6]_net_1\);
    
    \S[25]\ : AXOI3
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(2), C
         => alu_sel_coeff(0), Y => \S[25]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \S[17]\ : AO16
      port map(A => alu_sel_coeff(2), B => alu_sel_coeff(1), C
         => alu_sel_coeff(0), Y => \S[17]_net_1\);
    
    \S[10]\ : AO17
      port map(A => alu_sel_coeff(0), B => alu_sel_coeff(2), C
         => alu_sel_coeff(1), Y => \S[10]_net_1\);
    
    \S[20]\ : OA1A
      port map(A => alu_sel_coeff(2), B => alu_sel_coeff(0), C
         => alu_sel_coeff(1), Y => \S[20]_net_1\);
    
    \S[7]\ : AO16
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(0), C
         => alu_sel_coeff(2), Y => \S[7]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \S[18]\ : XAI1A
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff_0_2, C
         => alu_sel_coeff(1), Y => \S[19]\);
    
    \S[0]\ : AXO5
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff_0_2, C
         => alu_sel_coeff_0_0, Y => \S[0]_net_1\);
    
    \S[29]\ : OR3
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff(1), C
         => alu_sel_coeff_0_2, Y => \S[33]\);
    
    \S[1]\ : XNOR2
      port map(A => alu_sel_coeff_0_2, B => alu_sel_coeff_0_0, Y
         => \S_i[1]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \S[12]\ : AO1A
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff(1), C
         => alu_sel_coeff(2), Y => \S[12]_net_1\);
    
    \S[22]\ : AXO5
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff_0_2, C
         => alu_sel_coeff(1), Y => \S[22]_net_1\);
    
    \S[2]\ : NOR3B
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(2), C
         => alu_sel_coeff(0), Y => \S[2]_net_1\);
    
    \S[16]\ : MX2B
      port map(A => alu_sel_coeff_0_2, B => alu_sel_coeff_0_0, S
         => alu_sel_coeff(1), Y => \S[16]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MUXN_9_4 is

    port( alu_coef_s        : out   std_logic_vector(8 downto 0);
          S_0               : out   std_logic;
          S_i_0             : out   std_logic_vector(33 to 33);
          alu_sel_coeff     : in    std_logic_vector(4 downto 0);
          alu_sel_coeff_0_2 : in    std_logic;
          alu_sel_coeff_0_0 : in    std_logic
        );

end MUXN_9_4;

architecture DEF_ARCH of MUXN_9_4 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUXN_9_3
    port( alu_coef_s        : out   std_logic_vector(8 downto 0);
          S_0_0             : in    std_logic := 'U';
          S_0_18            : in    std_logic := 'U';
          alu_sel_coeff_0_0 : in    std_logic := 'U';
          alu_sel_coeff_0_2 : in    std_logic := 'U';
          alu_sel_coeff     : in    std_logic_vector(4 downto 0) := (others => 'U')
        );
  end component;

    signal \S[26]\, \S[8]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : MUXN_9_3
	Use entity work.MUXN_9_3(DEF_ARCH);
begin 

    S_0 <= \S[8]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \S[20]\ : OR2B
      port map(A => alu_sel_coeff(1), B => alu_sel_coeff(0), Y
         => \S[8]\);
    
    \S[18]\ : XOR2
      port map(A => alu_sel_coeff(0), B => alu_sel_coeff(1), Y
         => S_i_0(33));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \S[23]\ : NOR2A
      port map(A => alu_sel_coeff_0_0, B => alu_sel_coeff(1), Y
         => \S[26]\);
    
    \NB_STAGE_PLUS.MUXN_1\ : MUXN_9_3
      port map(alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0), S_0_0 => 
        \S[8]\, S_0_18 => \S[26]\, alu_sel_coeff_0_0 => 
        alu_sel_coeff_0_0, alu_sel_coeff_0_2 => alu_sel_coeff_0_2, 
        alu_sel_coeff(4) => alu_sel_coeff(4), alu_sel_coeff(3)
         => alu_sel_coeff(3), alu_sel_coeff(2) => 
        alu_sel_coeff(2), alu_sel_coeff(1) => alu_sel_coeff(1), 
        alu_sel_coeff(0) => alu_sel_coeff(0));
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MUXN_9_5 is

    port( alu_sel_coeff_0_0 : in    std_logic;
          alu_sel_coeff_0_2 : in    std_logic;
          alu_sel_coeff     : in    std_logic_vector(4 downto 0);
          S_i_0             : out   std_logic_vector(33 to 33);
          S                 : out   std_logic_vector(8 to 8);
          alu_coef_s        : out   std_logic_vector(8 downto 0)
        );

end MUXN_9_5;

architecture DEF_ARCH of MUXN_9_5 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MUXN_9_4
    port( alu_coef_s        : out   std_logic_vector(8 downto 0);
          S_0               : out   std_logic;
          S_i_0             : out   std_logic_vector(33 to 33);
          alu_sel_coeff     : in    std_logic_vector(4 downto 0) := (others => 'U');
          alu_sel_coeff_0_2 : in    std_logic := 'U';
          alu_sel_coeff_0_0 : in    std_logic := 'U'
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : MUXN_9_4
	Use entity work.MUXN_9_4(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \NB_STAGE_PLUS.MUXN_1\ : MUXN_9_4
      port map(alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0), S_0 => 
        S(8), S_i_0(33) => S_i_0(33), alu_sel_coeff(4) => 
        alu_sel_coeff(4), alu_sel_coeff(3) => alu_sel_coeff(3), 
        alu_sel_coeff(2) => alu_sel_coeff(2), alu_sel_coeff(1)
         => alu_sel_coeff(1), alu_sel_coeff(0) => 
        alu_sel_coeff(0), alu_sel_coeff_0_2 => alu_sel_coeff_0_2, 
        alu_sel_coeff_0_0 => alu_sel_coeff_0_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_18 is

    port( alu_sample : in    std_logic_vector(17 downto 0);
          OP1_2C_D   : out   std_logic_vector(17 downto 0);
          HRESETn_c  : in    std_logic;
          HCLK_c     : in    std_logic
        );

end MAC_REG_18;

architecture DEF_ARCH of MAC_REG_18 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Q[6]\ : DFN1C0
      port map(D => alu_sample(6), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(6));
    
    \Q[13]\ : DFN1C0
      port map(D => alu_sample(13), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(13));
    
    \Q[14]\ : DFN1C0
      port map(D => alu_sample(14), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(14));
    
    \Q[15]\ : DFN1C0
      port map(D => alu_sample(15), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(15));
    
    \Q[11]\ : DFN1C0
      port map(D => alu_sample(11), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(11));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Q[2]\ : DFN1C0
      port map(D => alu_sample(2), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(2));
    
    \Q[4]\ : DFN1C0
      port map(D => alu_sample(4), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(4));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Q[17]\ : DFN1C0
      port map(D => alu_sample(17), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(17));
    
    \Q[10]\ : DFN1C0
      port map(D => alu_sample(10), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(10));
    
    GND_i : GND
      port map(Y => \GND\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q[3]\ : DFN1C0
      port map(D => alu_sample(3), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(3));
    
    \Q[7]\ : DFN1C0
      port map(D => alu_sample(7), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(7));
    
    \Q[12]\ : DFN1C0
      port map(D => alu_sample(12), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(12));
    
    \Q[8]\ : DFN1C0
      port map(D => alu_sample(8), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(8));
    
    \Q[1]\ : DFN1C0
      port map(D => alu_sample(1), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(1));
    
    \Q[0]\ : DFN1C0
      port map(D => alu_sample(0), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(0));
    
    \Q[9]\ : DFN1C0
      port map(D => alu_sample(9), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(9));
    
    \Q[5]\ : DFN1C0
      port map(D => alu_sample(5), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(5));
    
    \Q[16]\ : DFN1C0
      port map(D => alu_sample(16), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP1_2C_D(16));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_9 is

    port( alu_coef_s : in    std_logic_vector(8 downto 0);
          OP2_2C_D   : out   std_logic_vector(8 downto 0);
          HRESETn_c  : in    std_logic;
          HCLK_c     : in    std_logic
        );

end MAC_REG_9;

architecture DEF_ARCH of MAC_REG_9 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Q[5]\ : DFN1C0
      port map(D => alu_coef_s(5), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(5));
    
    \Q[3]\ : DFN1C0
      port map(D => alu_coef_s(3), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(3));
    
    \Q[8]\ : DFN1C0
      port map(D => alu_coef_s(8), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(8));
    
    \Q[7]\ : DFN1C0
      port map(D => alu_coef_s(7), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(7));
    
    \Q[1]\ : DFN1C0
      port map(D => alu_coef_s(1), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(1));
    
    \Q[2]\ : DFN1C0
      port map(D => alu_coef_s(2), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(2));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q[6]\ : DFN1C0
      port map(D => alu_coef_s(6), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(6));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Q[0]\ : DFN1C0
      port map(D => alu_coef_s(0), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(0));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Q[4]\ : DFN1C0
      port map(D => alu_coef_s(4), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => OP2_2C_D(4));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_1_4 is

    port( MACMUX2sel_D   : in    std_logic;
          HRESETn_c      : in    std_logic;
          HCLK_c         : in    std_logic;
          MACMUX2sel_D_D : out   std_logic
        );

end MAC_REG_1_4;

architecture DEF_ARCH of MAC_REG_1_4 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q[0]\ : DFN1C0
      port map(D => MACMUX2sel_D, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MACMUX2sel_D_D);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_CONTROLER is

    port( alu_ctrl   : in    std_logic_vector(1 downto 0);
          MACMUX2sel : out   std_logic;
          N_4        : out   std_logic;
          mult       : out   std_logic;
          mult_0     : out   std_logic
        );

end MAC_CONTROLER;

architecture DEF_ARCH of MAC_CONTROLER is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un1_mult_i : NOR2B
      port map(A => alu_ctrl(1), B => alu_ctrl(0), Y => N_4);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un2_mult_i_x2 : XOR2
      port map(A => alu_ctrl(1), B => alu_ctrl(0), Y => mult);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un2_mult_i_x2_0 : XOR2
      port map(A => alu_ctrl(1), B => alu_ctrl(0), Y => mult_0);
    
    un1_add_0_a2 : NOR2A
      port map(A => alu_ctrl(1), B => alu_ctrl(0), Y => 
        MACMUX2sel);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_MUX is

    port( OP1_2C_D      : in    std_logic_vector(17 downto 0);
          MULTout       : in    std_logic_vector(24 downto 0);
          ADDERinB      : out   std_logic_vector(24 downto 0);
          ADDERinA_i    : out   std_logic_vector(18 to 18);
          OP2_2C_D      : in    std_logic_vector(8 downto 0);
          ADDERout      : in    std_logic_vector(24 downto 0);
          ADDERinA_17   : out   std_logic;
          ADDERinA_24   : out   std_logic;
          ADDERinA_23   : out   std_logic;
          ADDERinA_22   : out   std_logic;
          ADDERinA_21   : out   std_logic;
          ADDERinA_20   : out   std_logic;
          ADDERinA_19   : out   std_logic;
          ADDERinA_16   : out   std_logic;
          ADDERinA_15   : out   std_logic;
          ADDERinA_14   : out   std_logic;
          ADDERinA_13   : out   std_logic;
          ADDERinA_12   : out   std_logic;
          ADDERinA_11   : out   std_logic;
          ADDERinA_10   : out   std_logic;
          ADDERinA_9    : out   std_logic;
          ADDERinA_8    : out   std_logic;
          ADDERinA_7    : out   std_logic;
          ADDERinA_6    : out   std_logic;
          ADDERinA_5    : out   std_logic;
          ADDERinA_4    : out   std_logic;
          ADDERinA_3    : out   std_logic;
          ADDERinA_2    : out   std_logic;
          ADDERinA_1    : out   std_logic;
          ADDERinA_0    : out   std_logic;
          MACMUXsel_D   : in    std_logic;
          MACMUXsel_D_1 : in    std_logic;
          MACMUXsel_D_0 : in    std_logic
        );

end MAC_MUX;

architecture DEF_ARCH of MAC_MUX is 

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \OUTA[24]\ : MX2C
      port map(A => ADDERout(24), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_24);
    
    \OUTB[3]\ : MX2
      port map(A => MULTout(3), B => OP1_2C_D(3), S => 
        MACMUXsel_D_1, Y => ADDERinB(3));
    
    \OUTB[9]\ : MX2
      port map(A => MULTout(9), B => OP1_2C_D(9), S => 
        MACMUXsel_D_1, Y => ADDERinB(9));
    
    \OUTA[0]\ : MX2
      port map(A => ADDERout(0), B => OP2_2C_D(0), S => 
        MACMUXsel_D_0, Y => ADDERinA_0);
    
    \OUTA[3]\ : MX2
      port map(A => ADDERout(3), B => OP2_2C_D(3), S => 
        MACMUXsel_D_0, Y => ADDERinA_3);
    
    \OUTB[11]\ : MX2
      port map(A => MULTout(11), B => OP1_2C_D(11), S => 
        MACMUXsel_D, Y => ADDERinB(11));
    
    \OUTB[23]\ : MX2
      port map(A => MULTout(23), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(23));
    
    \OUTB[12]\ : MX2
      port map(A => MULTout(12), B => OP1_2C_D(12), S => 
        MACMUXsel_D, Y => ADDERinB(12));
    
    \OUTB[20]\ : MX2
      port map(A => MULTout(20), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(20));
    
    \OUTB[19]\ : MX2
      port map(A => MULTout(19), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(19));
    
    \OUTA[13]\ : MX2
      port map(A => ADDERout(13), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_13);
    
    \OUTB[8]\ : MX2
      port map(A => MULTout(8), B => OP1_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinB(8));
    
    \OUTA[10]\ : MX2
      port map(A => ADDERout(10), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_10);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \OUTB[6]\ : MX2
      port map(A => MULTout(6), B => OP1_2C_D(6), S => 
        MACMUXsel_D_1, Y => ADDERinB(6));
    
    \OUTA[6]\ : MX2
      port map(A => ADDERout(6), B => OP2_2C_D(6), S => 
        MACMUXsel_D_0, Y => ADDERinA_6);
    
    \OUTB[24]\ : MX2
      port map(A => MULTout(24), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(24));
    
    \OUTA[14]\ : MX2C
      port map(A => ADDERout(14), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_14);
    
    \OUTB[2]\ : MX2
      port map(A => MULTout(2), B => OP1_2C_D(2), S => 
        MACMUXsel_D_1, Y => ADDERinB(2));
    
    \OUTB[13]\ : MX2
      port map(A => MULTout(13), B => OP1_2C_D(13), S => 
        MACMUXsel_D, Y => ADDERinB(13));
    
    \OUTB[10]\ : MX2
      port map(A => MULTout(10), B => OP1_2C_D(10), S => 
        MACMUXsel_D, Y => ADDERinB(10));
    
    \OUTA[9]\ : MX2
      port map(A => ADDERout(9), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_9);
    
    \OUTA[15]\ : MX2C
      port map(A => ADDERout(15), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_15);
    
    \OUTA[16]\ : MX2
      port map(A => ADDERout(16), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_16);
    
    \OUTA[7]\ : MX2
      port map(A => ADDERout(7), B => OP2_2C_D(7), S => 
        MACMUXsel_D_0, Y => ADDERinA_7);
    
    \OUTB[5]\ : MX2
      port map(A => MULTout(5), B => OP1_2C_D(5), S => 
        MACMUXsel_D_1, Y => ADDERinB(5));
    
    \OUTB[14]\ : MX2
      port map(A => MULTout(14), B => OP1_2C_D(14), S => 
        MACMUXsel_D, Y => ADDERinB(14));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \OUTA[18]\ : MX2C
      port map(A => ADDERout(18), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_i(18));
    
    \OUTB[4]\ : MX2
      port map(A => MULTout(4), B => OP1_2C_D(4), S => 
        MACMUXsel_D_1, Y => ADDERinB(4));
    
    \OUTB[15]\ : MX2
      port map(A => MULTout(15), B => OP1_2C_D(15), S => 
        MACMUXsel_D, Y => ADDERinB(15));
    
    \OUTB[16]\ : MX2
      port map(A => MULTout(16), B => OP1_2C_D(16), S => 
        MACMUXsel_D, Y => ADDERinB(16));
    
    \OUTA[21]\ : MX2
      port map(A => ADDERout(21), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_21);
    
    \OUTA[22]\ : MX2C
      port map(A => ADDERout(22), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_22);
    
    \OUTA[17]\ : MX2
      port map(A => ADDERout(17), B => OP2_2C_D(8), S => 
        MACMUXsel_D, Y => ADDERinA_17);
    
    \OUTB[18]\ : MX2
      port map(A => MULTout(18), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(18));
    
    \OUTA[4]\ : MX2
      port map(A => ADDERout(4), B => OP2_2C_D(4), S => 
        MACMUXsel_D_0, Y => ADDERinA_4);
    
    \OUTA[1]\ : MX2C
      port map(A => ADDERout(1), B => OP2_2C_D(1), S => 
        MACMUXsel_D_0, Y => ADDERinA_1);
    
    \OUTB[7]\ : MX2
      port map(A => MULTout(7), B => OP1_2C_D(7), S => 
        MACMUXsel_D_1, Y => ADDERinB(7));
    
    \OUTA[2]\ : MX2
      port map(A => ADDERout(2), B => OP2_2C_D(2), S => 
        MACMUXsel_D_0, Y => ADDERinA_2);
    
    \OUTA[23]\ : MX2
      port map(A => ADDERout(23), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_23);
    
    \OUTA[20]\ : MX2
      port map(A => ADDERout(20), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_20);
    
    \OUTB[17]\ : MX2
      port map(A => MULTout(17), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(17));
    
    \OUTB[21]\ : MX2
      port map(A => MULTout(21), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(21));
    
    \OUTA[8]\ : MX2
      port map(A => ADDERout(8), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_8);
    
    \OUTB[22]\ : MX2
      port map(A => MULTout(22), B => OP1_2C_D(17), S => 
        MACMUXsel_D, Y => ADDERinB(22));
    
    \OUTB[0]\ : MX2
      port map(A => MULTout(0), B => OP1_2C_D(0), S => 
        MACMUXsel_D_1, Y => ADDERinB(0));
    
    \OUTA[11]\ : MX2
      port map(A => ADDERout(11), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_11);
    
    \OUTB[1]\ : MX2
      port map(A => MULTout(1), B => OP1_2C_D(1), S => 
        MACMUXsel_D_1, Y => ADDERinB(1));
    
    \OUTA[5]\ : MX2
      port map(A => ADDERout(5), B => OP2_2C_D(5), S => 
        MACMUXsel_D_0, Y => ADDERinA_5);
    
    \OUTA[12]\ : MX2
      port map(A => ADDERout(12), B => OP2_2C_D(8), S => 
        MACMUXsel_D_0, Y => ADDERinA_12);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \OUTA[19]\ : MX2
      port map(A => ADDERout(19), B => OP2_2C_D(8), S => 
        MACMUXsel_D_1, Y => ADDERinA_19);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_27 is

    port( MULTout   : in    std_logic_vector(24 downto 7);
          MULTout_D : out   std_logic_vector(24 downto 7);
          HRESETn_c : in    std_logic;
          HCLK_c    : in    std_logic
        );

end MAC_REG_27;

architecture DEF_ARCH of MAC_REG_27 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Q[24]\ : DFN1C0
      port map(D => MULTout(24), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(24));
    
    \Q[21]\ : DFN1C0
      port map(D => MULTout(21), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(21));
    
    \Q[13]\ : DFN1C0
      port map(D => MULTout(13), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(13));
    
    \Q[14]\ : DFN1C0
      port map(D => MULTout(14), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(14));
    
    \Q[15]\ : DFN1C0
      port map(D => MULTout(15), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(15));
    
    \Q[11]\ : DFN1C0
      port map(D => MULTout(11), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(11));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Q[20]\ : DFN1C0
      port map(D => MULTout(20), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(20));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Q[17]\ : DFN1C0
      port map(D => MULTout(17), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(17));
    
    \Q[10]\ : DFN1C0
      port map(D => MULTout(10), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(10));
    
    \Q[19]\ : DFN1C0
      port map(D => MULTout(19), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(19));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Q[18]\ : DFN1C0
      port map(D => MULTout(18), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(18));
    
    \Q[22]\ : DFN1C0
      port map(D => MULTout(22), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(22));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q[7]\ : DFN1C0
      port map(D => MULTout(7), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(7));
    
    \Q[12]\ : DFN1C0
      port map(D => MULTout(12), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(12));
    
    \Q[8]\ : DFN1C0
      port map(D => MULTout(8), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(8));
    
    \Q[9]\ : DFN1C0
      port map(D => MULTout(9), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(9));
    
    \Q[23]\ : DFN1C0
      port map(D => MULTout(23), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(23));
    
    \Q[16]\ : DFN1C0
      port map(D => MULTout(16), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MULTout_D(16));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_1_1 is

    port( alu_ctrl  : in    std_logic_vector(0 to 0);
          add_D     : out   std_logic;
          HRESETn_c : in    std_logic;
          HCLK_c    : in    std_logic;
          add_D_0   : out   std_logic
        );

end MAC_REG_1_1;

architecture DEF_ARCH of MAC_REG_1_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q_0[0]\ : DFN1C0
      port map(D => alu_ctrl(0), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => add_D_0);
    
    \Q[0]\ : DFN1C0
      port map(D => alu_ctrl(0), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => add_D);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_1_3 is

    port( MACMUX2sel   : in    std_logic;
          HRESETn_c    : in    std_logic;
          HCLK_c       : in    std_logic;
          MACMUX2sel_D : out   std_logic
        );

end MAC_REG_1_3;

architecture DEF_ARCH of MAC_REG_1_3 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q[0]\ : DFN1C0
      port map(D => MACMUX2sel, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => MACMUX2sel_D);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_1 is

    port( alu_ctrl    : in    std_logic_vector(2 to 2);
          clr_MAC_D   : out   std_logic;
          HRESETn_c   : in    std_logic;
          HCLK_c      : in    std_logic;
          clr_MAC_D_0 : out   std_logic
        );

end MAC_REG_1;

architecture DEF_ARCH of MAC_REG_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q_0[0]\ : DFN1C0
      port map(D => alu_ctrl(2), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => clr_MAC_D_0);
    
    \Q[0]\ : DFN1C0
      port map(D => alu_ctrl(2), CLK => HCLK_c, CLR => HRESETn_c, 
        Q => clr_MAC_D);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Adder is

    port( ADDERout     : out   std_logic_vector(24 downto 0);
          ADDERinA_i   : in    std_logic_vector(18 to 18);
          ADDERinB     : in    std_logic_vector(24 downto 0);
          ADDERinA_0   : in    std_logic;
          ADDERinA_1   : in    std_logic;
          ADDERinA_3   : in    std_logic;
          ADDERinA_5   : in    std_logic;
          ADDERinA_7   : in    std_logic;
          ADDERinA_8   : in    std_logic;
          ADDERinA_15  : in    std_logic;
          ADDERinA_16  : in    std_logic;
          ADDERinA_2   : in    std_logic;
          ADDERinA_14  : in    std_logic;
          ADDERinA_6   : in    std_logic;
          ADDERinA_10  : in    std_logic;
          ADDERinA_4   : in    std_logic;
          ADDERinA_12  : in    std_logic;
          ADDERinA_20  : in    std_logic;
          ADDERinA_11  : in    std_logic;
          ADDERinA_19  : in    std_logic;
          ADDERinA_9   : in    std_logic;
          ADDERinA_13  : in    std_logic;
          ADDERinA_21  : in    std_logic;
          ADDERinA_22  : in    std_logic;
          ADDERinA_24  : in    std_logic;
          ADDERinA_23  : in    std_logic;
          ADDERinA_17  : in    std_logic;
          HRESETn_c    : in    std_logic;
          HCLK_c       : in    std_logic;
          clr_MAC_D    : in    std_logic;
          add_D        : in    std_logic;
          clr_MAC_D_0  : in    std_logic;
          MACMUX2sel_D : in    std_logic;
          add_D_0      : in    std_logic
        );

end Adder;

architecture DEF_ARCH of Adder is 

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \un1_clr_1_0\, ADD_27x27_fast_I247_Y_0_0, 
        ADD_27x27_fast_I253_Y_0_0, ADD_27x27_fast_I254_Y_0_0, 
        ADD_27x27_fast_I208_Y_3, N534, N519, 
        ADD_27x27_fast_I208_Y_2, N472, N465, 
        ADD_27x27_fast_I208_Y_1, N415, N412, 
        ADD_27x27_fast_I208_Y_0, N388, ADD_27x27_fast_I251_Y_0_0, 
        ADD_27x27_fast_I207_Y_3, N532, N517, 
        ADD_27x27_fast_I207_Y_2, N470, N463, 
        ADD_27x27_fast_I207_Y_1, N413, N410, 
        ADD_27x27_fast_I207_Y_0, N391, ADD_27x27_fast_I243_Y_0_0, 
        ADD_27x27_fast_I239_Y_0_0, ADD_27x27_fast_I249_Y_0_0, 
        ADD_27x27_fast_I196_Y_0_0, N496, N_73, N439, 
        ADD_27x27_fast_I241_Y_0_0, ADD_27x27_fast_I250_Y_0_0, 
        ADD_27x27_fast_I242_Y_0_0, ADD_27x27_fast_I252_Y_0_0, 
        ADD_27x27_fast_I212_Y_1, N542, N527, 
        ADD_27x27_fast_I212_Y_0, N480, N473, 
        ADD_27x27_fast_I164_Y_i_0, N_58, 
        ADD_27x27_fast_I248_Y_0_0, ADD_27x27_fast_I211_Y_1, N540, 
        N525, ADD_27x27_fast_I211_Y_0, N478, N471, 
        ADD_27x27_fast_I209_Y_2, N536, N521, 
        ADD_27x27_fast_I209_Y_1, N474, N467, 
        ADD_27x27_fast_I209_Y_0, N417, N414, 
        ADD_27x27_fast_I240_Y_0_0, ADD_27x27_fast_I213_Y_1, 
        ADD_27x27_fast_I213_un1_Y_0, N529, 
        ADD_27x27_fast_I213_Y_0, N475, N482, 
        ADD_27x27_fast_I236_Y_0_0, N499, N_47, N491, 
        ADD_27x27_fast_I99_Y_0, N364, ADD_27x27_fast_I91_Y_0, 
        N376, ADD_27x27_fast_I107_Y_0, N352, 
        ADD_27x27_fast_I115_Y_0, N340, 
        ADD_27x27_fast_I115_un1_Y_0, N_108, 
        ADD_27x27_fast_I116_Y_0, ADD_27x27_fast_I100_Y_0, N362, 
        I207_un1_Y, N533, N548, I209_un1_Y, N537, N552, 
        I211_un1_Y, N541, N502, N431, N428, N481, N488, N436, 
        N444, N497, I208_un1_Y, N535, N550, I212_un1_Y, N543, 
        N_48, N_33, \un1_clr_1\, \un2_resadd[24]\, 
        \un2_resadd[23]\, \un2_resadd[22]\, \un2_resadd[21]\, 
        ADD_27x27_fast_I210_Y_0_a2, \un2_resadd[20]\, 
        \un2_resadd[19]\, \un2_resadd[18]\, I185_un1_Y, 
        \un2_resadd[16]\, N648_i, \un2_resadd[15]\, N651, 
        \un2_resadd[14]\, N654_i, \un2_resadd[13]\, 
        ADD_27x27_fast_I192_Y_0_a2, N361, \un2_resadd[12]\, 
        I193_un1_Y, \un2_resadd[11]\, I194_un1_Y_i, 
        \un2_resadd[10]\, N544, I195_un1_Y_i, \un2_resadd[9]\, 
        N_78_i, \un2_resadd[8]\, \un2_resadd[7]\, \un2_resadd[6]\, 
        \un2_resadd[5]\, \un2_resadd[4]\, \un2_resadd[3]\, 
        \un2_resadd[2]\, \un2_resadd[1]\, N325, \un2_resadd[17]\, 
        N423, N_98_i, N420, N392, N355, N356, N379, N380, N385, 
        N386, N429, N437, N349, N441, N343, N445, N_52_i_0, N449, 
        N_72, N450, N418, N433, N430, N483, N434, N490, N438, 
        N442, N494, N498, N446, N487, N479, N495, I163_un1_Y, 
        N383, N350, N344, N341, N486, N346, N382, N367, N368, 
        N_105_1, N489, I190_un1_Y, N_59, N_50, N_9, N_11, N_16, 
        N_18, N_23, N_30, N_32, \REG_4[1]\, \REG_4[3]\, 
        \REG_4[8]\, \REG_4[10]\, \REG_4[15]\, \REG_4[22]\, 
        \REG_4[24]\, N_8, N_12, N_15, N_19, N_22, N_26, N_29, 
        \REG_4[0]\, \REG_4[4]\, \REG_4[7]\, \REG_4[11]\, 
        \REG_4[14]\, \REG_4[18]\, \REG_4[21]\, N_10, N_13, N_14, 
        N_17, N_20, N_21, N_24, N_27, N_28, N_31, \REG_4[2]\, 
        \REG_4[5]\, \REG_4[6]\, \REG_4[9]\, \REG_4[12]\, 
        \REG_4[13]\, \REG_4[16]\, \REG_4[19]\, \REG_4[20]\, 
        \REG_4[23]\, N_23_0, \REG_4[17]\, N_25, N374, N370, N373, 
        N371, N426, N422, N421, N425, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    un2_resadd_ADD_27x27_fast_I8_G0N : NOR2B
      port map(A => ADDERinB(8), B => ADDERinA_8, Y => N349);
    
    un2_resadd_ADD_27x27_fast_I241_Y_0_0 : XOR2
      port map(A => ADDERinA_11, B => ADDERinB(11), Y => 
        ADD_27x27_fast_I241_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I134_Y : NOR2
      port map(A => N475, B => N467, Y => N521);
    
    un2_resadd_ADD_27x27_fast_I208_Y_1 : AOI1B
      port map(A => N415, B => N412, C => ADD_27x27_fast_I208_Y_0, 
        Y => ADD_27x27_fast_I208_Y_1);
    
    un2_resadd_ADD_27x27_fast_I156_Y : NOR2A
      port map(A => N497, B => N489, Y => N543);
    
    un2_resadd_ADD_27x27_fast_I19_P0N : OR2
      port map(A => ADDERinB(19), B => ADDERinA_19, Y => N383);
    
    un2_resadd_ADD_27x27_fast_I21_G0N : NOR2B
      port map(A => ADDERinB(21), B => ADDERinA_21, Y => N388);
    
    \REG[14]\ : DFN1E0C0
      port map(D => \REG_4[14]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(14));
    
    un2_resadd_ADD_27x27_fast_I214_Y_0_a2 : OR2A
      port map(A => N651, B => N_23_0, Y => N_98_i);
    
    un2_resadd_ADD_27x27_fast_I12_G0N : OR2B
      port map(A => ADDERinB(12), B => ADDERinA_12, Y => N361);
    
    un2_resadd_ADD_27x27_fast_I99_Y : AOI1
      port map(A => N431, B => N428, C => ADD_27x27_fast_I99_Y_0, 
        Y => N480);
    
    un2_resadd_ADD_27x27_fast_I149_Y : AO1A
      port map(A => N483, B => N490, C => N482, Y => N536);
    
    un2_resadd_ADD_27x27_fast_I68_Y : OA1
      port map(A => ADDERinA_4, B => ADDERinB(4), C => N341, Y
         => N446);
    
    un2_resadd_ADD_27x27_fast_I5_P0N : OR2
      port map(A => ADDERinB(5), B => ADDERinA_5, Y => N341);
    
    un2_resadd_ADD_27x27_fast_I11_G0N_0_o2 : OR2B
      port map(A => ADDERinB(11), B => ADDERinA_11, Y => N_50);
    
    un2_resadd_ADD_27x27_fast_I209_Y_0 : AOI1
      port map(A => N417, B => N414, C => N413, Y => 
        ADD_27x27_fast_I209_Y_0);
    
    un2_resadd_ADD_27x27_fast_I132_Y : NOR2
      port map(A => N473, B => N465, Y => N519);
    
    un2_resadd_ADD_27x27_fast_I122_Y_i_o2 : MAJ3
      port map(A => ADDERinA_2, B => ADDERinB(2), C => N_47, Y
         => N_48);
    
    un2_resadd_ADD_27x27_fast_I93_Y : AO1
      port map(A => N425, B => N422, C => N421, Y => N474);
    
    un2_resadd_ADD_27x27_fast_I52_Y : OA1
      port map(A => ADDERinA_13, B => ADDERinB(13), C => N362, Y
         => N430);
    
    un2_resadd_ADD_27x27_fast_I254_Y_0 : AX1C
      port map(A => I207_un1_Y, B => ADD_27x27_fast_I207_Y_3, C
         => ADD_27x27_fast_I254_Y_0_0, Y => \un2_resadd[24]\);
    
    \REG_RNO[11]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_19, Y => \REG_4[11]\);
    
    \REG[22]\ : DFN1E0C0
      port map(D => \REG_4[22]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(22));
    
    un2_resadd_ADD_27x27_fast_I51_Y : AO13
      port map(A => ADDERinB(13), B => ADDERinA_13, C => N361, Y
         => N429);
    
    \REG_RNO[20]\ : NOR2
      port map(A => clr_MAC_D, B => N_28, Y => \REG_4[20]\);
    
    \REG_RNO[15]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_23, Y => \REG_4[15]\);
    
    \REG_RNO_0[17]\ : MX2C
      port map(A => ADDERinB(17), B => \un2_resadd[17]\, S => 
        add_D, Y => N_25);
    
    un2_resadd_ADD_27x27_fast_I196_Y_0_a2 : OR3B
      port map(A => N497, B => N_48, C => N_73, Y => N_78_i);
    
    un2_resadd_ADD_27x27_fast_I240_Y_0_0 : XOR2
      port map(A => ADDERinA_10, B => ADDERinB(10), Y => 
        ADD_27x27_fast_I240_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I6_G0N : NOR2B
      port map(A => ADDERinB(6), B => ADDERinA_6, Y => N343);
    
    un2_resadd_ADD_27x27_fast_I163_Y : OR2
      port map(A => N498, B => I163_un1_Y, Y => N552);
    
    un2_resadd_ADD_27x27_fast_I90_Y : OR2B
      port map(A => N422, B => N418, Y => N471);
    
    un2_resadd_ADD_27x27_fast_I35_Y : MAJ3
      port map(A => ADDERinA_21, B => ADDERinB(21), C => N385, Y
         => N413);
    
    un2_resadd_ADD_27x27_fast_I48_Y : NOR2B
      port map(A => N371, B => N368, Y => N426);
    
    \REG_RNO[9]\ : NOR2
      port map(A => clr_MAC_D, B => N_17, Y => \REG_4[9]\);
    
    \REG_RNO_0[8]\ : MX2C
      port map(A => ADDERinB(8), B => \un2_resadd[8]\, S => 
        add_D_0, Y => N_16);
    
    \REG[11]\ : DFN1E0C0
      port map(D => \REG_4[11]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(11));
    
    un2_resadd_ADD_27x27_fast_I99_Y_0 : AO18
      port map(A => N364, B => ADDERinB(14), C => ADDERinA_14, Y
         => ADD_27x27_fast_I99_Y_0);
    
    un2_resadd_ADD_27x27_fast_I6_P0N : OR2
      port map(A => ADDERinB(6), B => ADDERinA_6, Y => N344);
    
    un2_resadd_ADD_27x27_fast_I15_G0N : NOR2A
      port map(A => ADDERinB(15), B => ADDERinA_15, Y => N370);
    
    un2_resadd_ADD_27x27_fast_I207_Y_1 : AOI1B
      port map(A => N413, B => N410, C => ADD_27x27_fast_I207_Y_0, 
        Y => ADD_27x27_fast_I207_Y_1);
    
    un2_resadd_ADD_27x27_fast_I207_Y_0 : MIN3
      port map(A => ADDERinA_23, B => ADDERinB(23), C => N391, Y
         => ADD_27x27_fast_I207_Y_0);
    
    un2_resadd_ADD_27x27_fast_I116_Y : NOR2B
      port map(A => ADD_27x27_fast_I116_Y_0, B => N444, Y => N497);
    
    un2_resadd_ADD_27x27_fast_I242_Y_0_0 : XOR2
      port map(A => ADDERinA_12, B => ADDERinB(12), Y => 
        ADD_27x27_fast_I242_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I163_un1_Y : NOR2B
      port map(A => N_47, B => N499, Y => I163_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I238_Y_0 : XOR3
      port map(A => ADDERinB(8), B => ADDERinA_8, C => N548, Y
         => \un2_resadd[8]\);
    
    \REG_RNO[4]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_12, Y => \REG_4[4]\);
    
    \REG_RNO[12]\ : NOR2
      port map(A => clr_MAC_D, B => N_20, Y => \REG_4[12]\);
    
    un2_resadd_ADD_27x27_fast_I140_Y : NOR2
      port map(A => N481, B => N473, Y => N527);
    
    un2_resadd_ADD_27x27_fast_I248_Y_0 : AX1B
      port map(A => I185_un1_Y, B => ADD_27x27_fast_I213_Y_1, C
         => ADD_27x27_fast_I248_Y_0_0, Y => \un2_resadd[18]\);
    
    \REG_RNO_0[11]\ : MX2C
      port map(A => ADDERinB(11), B => \un2_resadd[11]\, S => 
        add_D_0, Y => N_19);
    
    un2_resadd_ADD_27x27_fast_I66_Y : NOR2B
      port map(A => N344, B => N341, Y => N444);
    
    un2_resadd_ADD_27x27_fast_I247_Y_0_0 : XOR2
      port map(A => ADDERinA_17, B => ADDERinB(17), Y => 
        ADD_27x27_fast_I247_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I162_Y : AO1
      port map(A => N_48, B => N497, C => N496, Y => N550);
    
    un2_resadd_ADD_27x27_fast_I36_Y : OA1
      port map(A => ADDERinA_21, B => ADDERinB(21), C => N386, Y
         => N414);
    
    un2_resadd_ADD_27x27_fast_I209_Y_2 : AOI1B
      port map(A => N536, B => N521, C => ADD_27x27_fast_I209_Y_1, 
        Y => ADD_27x27_fast_I209_Y_2);
    
    un2_resadd_ADD_27x27_fast_I236_Y_0_0 : XOR2
      port map(A => ADDERinA_6, B => ADDERinB(6), Y => 
        ADD_27x27_fast_I236_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I212_Y_1 : AO1
      port map(A => N542, B => N527, C => ADD_27x27_fast_I212_Y_0, 
        Y => ADD_27x27_fast_I212_Y_1);
    
    un2_resadd_ADD_27x27_fast_I19_G0N : NOR2B
      port map(A => ADDERinB(19), B => ADDERinA_19, Y => N382);
    
    \REG_RNO_0[10]\ : MX2C
      port map(A => ADDERinB(10), B => \un2_resadd[10]\, S => 
        add_D_0, Y => N_18);
    
    \REG[12]\ : DFN1E0C0
      port map(D => \REG_4[12]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(12));
    
    un2_resadd_ADD_27x27_fast_I84_Y : OR2B
      port map(A => N_105_1, B => N412, Y => N465);
    
    un2_resadd_ADD_27x27_fast_I107_Y_0 : MIN3
      port map(A => ADDERinA_10, B => ADDERinB(10), C => N352, Y
         => ADD_27x27_fast_I107_Y_0);
    
    un2_resadd_ADD_27x27_fast_I185_un1_Y : NOR2B
      port map(A => N544, B => N529, Y => I185_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I115_un1_Y_0 : OA1B
      port map(A => ADDERinA_4, B => ADDERinB(4), C => N_108, Y
         => ADD_27x27_fast_I115_un1_Y_0);
    
    un2_resadd_ADD_27x27_fast_I207_Y_2 : OA1A
      port map(A => N470, B => N463, C => ADD_27x27_fast_I207_Y_1, 
        Y => ADD_27x27_fast_I207_Y_2);
    
    un2_resadd_ADD_27x27_fast_I118_Y : NOR2B
      port map(A => N450, B => N446, Y => N499);
    
    un2_resadd_ADD_27x27_fast_I207_Y_3 : AOI1B
      port map(A => N532, B => N517, C => ADD_27x27_fast_I207_Y_2, 
        Y => ADD_27x27_fast_I207_Y_3);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \REG_RNO_0[21]\ : MX2C
      port map(A => ADDERinB(21), B => \un2_resadd[21]\, S => 
        add_D, Y => N_29);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un2_resadd_ADD_27x27_fast_I63_Y : MAJ3
      port map(A => ADDERinA_7, B => ADDERinB(7), C => N343, Y
         => N441);
    
    un2_resadd_ADD_27x27_fast_I236_Y_0 : XOR2
      port map(A => ADD_27x27_fast_I236_Y_0_0, B => N552, Y => 
        \un2_resadd[6]\);
    
    un2_resadd_ADD_27x27_fast_I45_Y_0_o2 : AO1
      port map(A => N374, B => N370, C => N373, Y => N423);
    
    un2_resadd_ADD_27x27_fast_I10_G0N : NOR2B
      port map(A => ADDERinB(10), B => ADDERinA_10, Y => N355);
    
    un2_resadd_ADD_27x27_fast_I246_Y_0 : XNOR3
      port map(A => ADDERinB(16), B => ADDERinA_16, C => N648_i, 
        Y => \un2_resadd[16]\);
    
    \REG_RNO[14]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_22, Y => \REG_4[14]\);
    
    un2_resadd_ADD_27x27_fast_I92_Y : OR2A
      port map(A => N420, B => N_23_0, Y => N473);
    
    un2_resadd_ADD_27x27_fast_I39_Y : MAJ3
      port map(A => ADDERinA_19, B => ADDERinB(19), C => N379, Y
         => N417);
    
    un2_resadd_ADD_27x27_fast_I150_Y : NOR2
      port map(A => N491, B => N483, Y => N537);
    
    un2_resadd_ADD_27x27_fast_I235_Y_0 : XNOR3
      port map(A => ADDERinB(5), B => ADDERinA_5, C => N_33, Y
         => \un2_resadd[5]\);
    
    un2_resadd_ADD_27x27_fast_I164_Y_i_0 : MAJ3
      port map(A => ADDERinA_4, B => ADDERinB(4), C => N_58, Y
         => ADD_27x27_fast_I164_Y_i_0);
    
    un2_resadd_ADD_27x27_fast_I212_Y_0 : AO1D
      port map(A => N480, B => N473, C => N472, Y => 
        ADD_27x27_fast_I212_Y_0);
    
    un2_resadd_ADD_27x27_fast_I196_Y_0_0 : OA1C
      port map(A => N496, B => N_73, C => N439, Y => 
        ADD_27x27_fast_I196_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I245_Y_0 : XNOR3
      port map(A => ADDERinB(15), B => ADDERinA_15, C => N651, Y
         => \un2_resadd[15]\);
    
    \REG[0]\ : DFN1E0C0
      port map(D => \REG_4[0]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(0));
    
    \REG_RNO[7]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_15, Y => \REG_4[7]\);
    
    un2_resadd_ADD_27x27_fast_I9_G0N : NOR2B
      port map(A => ADDERinB(9), B => ADDERinA_9, Y => N352);
    
    un2_resadd_ADD_27x27_fast_I91_Y : AO1
      port map(A => N423, B => N420, C => ADD_27x27_fast_I91_Y_0, 
        Y => N472);
    
    \REG_RNO_0[20]\ : MX2C
      port map(A => ADDERinB(20), B => \un2_resadd[20]\, S => 
        add_D, Y => N_28);
    
    un2_resadd_ADD_27x27_fast_I212_un1_Y : NOR3C
      port map(A => N543, B => N527, C => N_48, Y => I212_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I106_Y : OR2B
      port map(A => N438, B => N434, Y => N487);
    
    un2_resadd_ADD_27x27_fast_I3_G0N_i_o2 : NOR2B
      port map(A => ADDERinB(3), B => ADDERinA_3, Y => N_59);
    
    un2_resadd_ADD_27x27_fast_I60_Y : OA1
      port map(A => ADDERinA_9, B => ADDERinB(9), C => N350, Y
         => N438);
    
    \REG[23]\ : DFN1E0C0
      port map(D => \REG_4[23]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(23));
    
    un2_resadd_ADD_27x27_fast_I208_Y_0 : AO18
      port map(A => N388, B => ADDERinA_22, C => ADDERinB(22), Y
         => ADD_27x27_fast_I208_Y_0);
    
    \REG_RNO[1]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_9, Y => \REG_4[1]\);
    
    un2_resadd_ADD_27x27_fast_I43_Y : MAJ3
      port map(A => ADDERinA_17, B => ADDERinB(17), C => N373, Y
         => N421);
    
    un2_resadd_ADD_27x27_fast_I190_un1_Y : NOR2B
      port map(A => N550, B => N535, Y => I190_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I20_P0N : OR2
      port map(A => ADDERinB(20), B => ADDERinA_20, Y => N386);
    
    un2_resadd_ADD_27x27_fast_I208_Y_2 : OA1A
      port map(A => N472, B => N465, C => ADD_27x27_fast_I208_Y_1, 
        Y => ADD_27x27_fast_I208_Y_2);
    
    un2_resadd_ADD_27x27_fast_I101_Y : AO1
      port map(A => N433, B => N430, C => N429, Y => N482);
    
    \REG_RNO[21]\ : NOR2
      port map(A => clr_MAC_D, B => N_29, Y => \REG_4[21]\);
    
    un2_resadd_ADD_27x27_fast_I16_G0N : NOR2B
      port map(A => ADDERinB(16), B => ADDERinA_16, Y => N373);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un2_resadd_ADD_27x27_fast_I91_Y_0 : AO13
      port map(A => N376, B => ADDERinB(18), C => ADDERinA_i(18), 
        Y => ADD_27x27_fast_I91_Y_0);
    
    un2_resadd_ADD_27x27_fast_I211_Y_0 : OA1C
      port map(A => N478, B => N471, C => N470, Y => 
        ADD_27x27_fast_I211_Y_0);
    
    un2_resadd_ADD_27x27_fast_I97_Y : AO1
      port map(A => N429, B => N426, C => N425, Y => N478);
    
    un2_resadd_ADD_27x27_fast_I40_Y : NOR2B
      port map(A => N383, B => N380, Y => N418);
    
    un2_resadd_ADD_27x27_fast_I2_G0N_i_o2 : OR2B
      port map(A => ADDERinB(2), B => ADDERinA_2, Y => N_72);
    
    \REG_RNO[13]\ : NOR2
      port map(A => clr_MAC_D, B => N_21, Y => \REG_4[13]\);
    
    un2_resadd_ADD_27x27_fast_I145_Y : AO1A
      port map(A => N479, B => N486, C => N478, Y => N532);
    
    un2_resadd_ADD_27x27_fast_I108_Y : OR2A
      port map(A => N436, B => N_73, Y => N489);
    
    \REG_RNO_0[19]\ : MX2C
      port map(A => ADDERinB(19), B => \un2_resadd[19]\, S => 
        add_D, Y => N_27);
    
    un2_resadd_ADD_27x27_fast_I110_Y : OR2B
      port map(A => N442, B => N438, Y => N491);
    
    \REG_RNO_0[6]\ : MX2C
      port map(A => ADDERinB(6), B => \un2_resadd[6]\, S => add_D, 
        Y => N_14);
    
    un2_resadd_ADD_27x27_fast_I22_P0N : OR2A
      port map(A => ADDERinA_22, B => ADDERinB(22), Y => N392);
    
    un2_resadd_ADD_27x27_fast_I213_Y_1 : AO1
      port map(A => ADD_27x27_fast_I213_un1_Y_0, B => N529, C => 
        ADD_27x27_fast_I213_Y_0, Y => ADD_27x27_fast_I213_Y_1);
    
    un2_resadd_ADD_27x27_fast_I72_Y : OA1
      port map(A => ADDERinA_2, B => ADDERinB(2), C => N_58, Y
         => N450);
    
    un2_resadd_ADD_27x27_fast_I116_Y_0 : OA1
      port map(A => ADDERinA_4, B => ADDERinB(4), C => N_58, Y
         => ADD_27x27_fast_I116_Y_0);
    
    un2_resadd_ADD_27x27_fast_I109_Y : AO1
      port map(A => N441, B => N438, C => N437, Y => N490);
    
    \REG[9]\ : DFN1E0C0
      port map(D => \REG_4[9]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(9));
    
    un1_clr_1_0 : NOR3
      port map(A => add_D_0, B => MACMUX2sel_D, C => clr_MAC_D_0, 
        Y => \un1_clr_1_0\);
    
    un2_resadd_ADD_27x27_fast_I142_Y : NOR2
      port map(A => N483, B => N475, Y => N529);
    
    \REG_RNO_0[9]\ : MX2C
      port map(A => ADDERinB(9), B => \un2_resadd[9]\, S => add_D, 
        Y => N_17);
    
    un2_resadd_ADD_27x27_fast_I71_Y : AO13
      port map(A => ADDERinB(3), B => ADDERinA_3, C => N_72, Y
         => N449);
    
    \REG_RNO[22]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_30, Y => \REG_4[22]\);
    
    \REG[5]\ : DFN1E0C0
      port map(D => \REG_4[5]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(5));
    
    un2_resadd_ADD_27x27_fast_I210_Y_0_a2 : OA1
      port map(A => I212_un1_Y, B => ADD_27x27_fast_I212_Y_1, C
         => N_105_1, Y => ADD_27x27_fast_I210_Y_0_a2);
    
    \REG_RNO[2]\ : NOR2
      port map(A => clr_MAC_D, B => N_10, Y => \REG_4[2]\);
    
    \REG[13]\ : DFN1E0C0
      port map(D => \REG_4[13]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(13));
    
    un2_resadd_ADD_27x27_fast_I153_Y : AO1A
      port map(A => N487, B => N494, C => N486, Y => N540);
    
    un2_resadd_ADD_27x27_fast_I232_Y_0 : XOR3
      port map(A => ADDERinB(2), B => ADDERinA_2, C => N_47, Y
         => \un2_resadd[2]\);
    
    un2_resadd_ADD_27x27_fast_I100_Y_0 : OA1
      port map(A => ADDERinA_11, B => ADDERinB(11), C => N362, Y
         => ADD_27x27_fast_I100_Y_0);
    
    \REG[6]\ : DFN1E0C0
      port map(D => \REG_4[6]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(6));
    
    \REG[18]\ : DFN1E0C0
      port map(D => \REG_4[18]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(18));
    
    un2_resadd_ADD_27x27_fast_I8_P0N : OR2
      port map(A => ADDERinB(8), B => ADDERinA_8, Y => N350);
    
    un2_resadd_ADD_27x27_fast_I14_G0N : NOR2A
      port map(A => ADDERinB(14), B => ADDERinA_14, Y => N367);
    
    un2_resadd_ADD_27x27_fast_I242_Y_0 : AX1D
      port map(A => I193_un1_Y, B => N540, C => 
        ADD_27x27_fast_I242_Y_0_0, Y => \un2_resadd[12]\);
    
    un2_resadd_ADD_27x27_fast_I211_un1_Y : OR3C
      port map(A => N525, B => N541, C => N502, Y => I211_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I46_Y_i : OR2B
      port map(A => N374, B => N371, Y => N_23_0);
    
    un2_resadd_ADD_27x27_fast_I239_Y_0_0 : XOR2
      port map(A => ADDERinA_9, B => ADDERinB(9), Y => 
        ADD_27x27_fast_I239_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I155_Y : AO1A
      port map(A => N489, B => N496, C => N488, Y => N542);
    
    un2_resadd_ADD_27x27_fast_I191_Y : AOI1
      port map(A => N552, B => N537, C => N536, Y => N654_i);
    
    \REG_RNO_0[13]\ : MX2C
      port map(A => ADDERinB(13), B => \un2_resadd[13]\, S => 
        add_D, Y => N_21);
    
    un2_resadd_ADD_27x27_fast_I249_Y_0_0 : XOR2
      port map(A => ADDERinA_19, B => ADDERinB(19), Y => 
        ADD_27x27_fast_I249_Y_0_0);
    
    \REG_RNO_0[18]\ : MX2C
      port map(A => ADDERinB(18), B => \un2_resadd[18]\, S => 
        add_D, Y => N_26);
    
    \REG_RNO[18]\ : NOR2
      port map(A => clr_MAC_D, B => N_26, Y => \REG_4[18]\);
    
    \REG[19]\ : DFN1E0C0
      port map(D => \REG_4[19]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(19));
    
    un2_resadd_ADD_27x27_fast_I32_Y : OA1
      port map(A => ADDERinA_23, B => ADDERinB(23), C => N392, Y
         => N410);
    
    un2_resadd_ADD_27x27_fast_I53_Y_0 : AO1C
      port map(A => N_50, B => N362, C => N361, Y => N431);
    
    un2_resadd_ADD_27x27_fast_I209_un1_Y : OR3C
      port map(A => N537, B => N521, C => N552, Y => I209_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I147_Y : AO1C
      port map(A => N481, B => N488, C => N480, Y => N534);
    
    un2_resadd_ADD_27x27_fast_I253_Y_0_0 : XOR2
      port map(A => ADDERinA_23, B => ADDERinB(23), Y => 
        ADD_27x27_fast_I253_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I7_G0N : NOR2B
      port map(A => ADDERinB(7), B => ADDERinA_7, Y => N346);
    
    un2_resadd_ADD_27x27_fast_I5_G0N : NOR2B
      port map(A => ADDERinB(5), B => ADDERinA_5, Y => N340);
    
    un2_resadd_ADD_27x27_fast_I138_Y : NOR2
      port map(A => N479, B => N471, Y => N525);
    
    un2_resadd_ADD_27x27_fast_I154_Y : NOR2A
      port map(A => N495, B => N487, Y => N541);
    
    un2_resadd_ADD_27x27_fast_I37_Y_0_o2 : AO1
      port map(A => N386, B => N382, C => N385, Y => N415);
    
    \REG_RNO[19]\ : NOR2
      port map(A => clr_MAC_D, B => N_27, Y => \REG_4[19]\);
    
    un2_resadd_ADD_27x27_fast_I58_Y : OA1
      port map(A => ADDERinA_9, B => ADDERinB(9), C => N356, Y
         => N436);
    
    \REG_RNO_0[1]\ : MX2C
      port map(A => ADDERinB(1), B => \un2_resadd[1]\, S => 
        add_D_0, Y => N_9);
    
    un2_resadd_ADD_27x27_fast_I94_Y : OR2B
      port map(A => N426, B => N422, Y => N475);
    
    un2_resadd_ADD_27x27_fast_I42_Y : OA1
      port map(A => ADDERinA_17, B => ADDERinB(17), C => N380, Y
         => N420);
    
    un2_resadd_ADD_27x27_fast_I86_Y : OR2B
      port map(A => N418, B => N414, Y => N467);
    
    un2_resadd_ADD_27x27_fast_I75_Y_i_o2 : AO18
      port map(A => ADDERinA_1, B => ADDERinB(1), C => N325, Y
         => N_47);
    
    un2_resadd_ADD_27x27_fast_I231_Y_0 : XOR3
      port map(A => ADDERinB(1), B => ADDERinA_1, C => N325, Y
         => \un2_resadd[1]\);
    
    \REG[1]\ : DFN1E0C0
      port map(D => \REG_4[1]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(1));
    
    un2_resadd_ADD_27x27_fast_I241_Y_0 : AX1A
      port map(A => N542, B => I194_un1_Y_i, C => 
        ADD_27x27_fast_I241_Y_0_0, Y => \un2_resadd[11]\);
    
    un2_resadd_ADD_27x27_fast_I17_G0N : NOR2B
      port map(A => ADDERinB(17), B => ADDERinA_17, Y => N376);
    
    un2_resadd_ADD_27x27_fast_I100_Y : OR2B
      port map(A => ADD_27x27_fast_I100_Y_0, B => N428, Y => N481);
    
    \REG_RNO[24]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_32, Y => \REG_4[24]\);
    
    un2_resadd_ADD_27x27_fast_I55_Y : MAJ3
      port map(A => ADDERinA_11, B => ADDERinB(11), C => N355, Y
         => N433);
    
    un2_resadd_ADD_27x27_fast_I193_un1_Y : NOR2B
      port map(A => N541, B => N502, Y => I193_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I164_Y_i : AO1C
      port map(A => N_48, B => N_108, C => 
        ADD_27x27_fast_I164_Y_i_0, Y => N_33);
    
    \REG[20]\ : DFN1E0C0
      port map(D => \REG_4[20]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(20));
    
    un2_resadd_ADD_27x27_fast_I252_Y_0 : AX1C
      port map(A => I209_un1_Y, B => ADD_27x27_fast_I209_Y_2, C
         => ADD_27x27_fast_I252_Y_0_0, Y => \un2_resadd[22]\);
    
    \REG_RNO[8]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_16, Y => \REG_4[8]\);
    
    \REG_RNO_0[7]\ : MX2C
      port map(A => ADDERinB(7), B => \un2_resadd[7]\, S => 
        add_D_0, Y => N_15);
    
    un2_resadd_ADD_27x27_fast_I67_Y : MAJ3
      port map(A => ADDERinA_5, B => ADDERinB(5), C => N_52_i_0, 
        Y => N445);
    
    \REG_RNO_0[23]\ : MX2C
      port map(A => ADDERinB(23), B => \un2_resadd[23]\, S => 
        add_D, Y => N_31);
    
    \REG[3]\ : DFN1E0C0
      port map(D => \REG_4[3]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(3));
    
    un2_resadd_ADD_27x27_fast_I248_Y_0_0 : XOR2
      port map(A => ADDERinA_i(18), B => ADDERinB(18), Y => 
        ADD_27x27_fast_I248_Y_0_0);
    
    \REG_RNO[3]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_11, Y => \REG_4[3]\);
    
    un2_resadd_ADD_27x27_fast_I121_Y : AO1
      port map(A => N_47, B => N450, C => N449, Y => N502);
    
    un2_resadd_ADD_27x27_fast_I113_Y : AO1
      port map(A => N445, B => N442, C => N441, Y => N494);
    
    \REG[17]\ : DFN1E0C0
      port map(D => \REG_4[17]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(17));
    
    un2_resadd_ADD_27x27_fast_I161_Y : AO1
      port map(A => N502, B => N495, C => N494, Y => N548);
    
    un2_resadd_ADD_27x27_fast_I22_G0N : NOR2A
      port map(A => ADDERinB(22), B => ADDERinA_22, Y => N391);
    
    un2_resadd_ADD_27x27_fast_I157_Y : AO1A
      port map(A => N491, B => N498, C => N490, Y => N544);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un2_resadd_ADD_27x27_fast_I195_un1_Y : OR3B
      port map(A => N499, B => N_47, C => N491, Y => I195_un1_Y_i);
    
    un2_resadd_ADD_27x27_fast_I115_Y : AO1B
      port map(A => ADD_27x27_fast_I115_un1_Y_0, B => N444, C => 
        ADD_27x27_fast_I115_Y_0, Y => N496);
    
    un2_resadd_ADD_27x27_fast_I89_Y : AO1
      port map(A => N421, B => N418, C => N417, Y => N470);
    
    \REG_RNO_0[16]\ : MX2C
      port map(A => ADDERinB(16), B => \un2_resadd[16]\, S => 
        add_D, Y => N_24);
    
    un2_resadd_ADD_27x27_fast_I213_Y_0 : AO1A
      port map(A => N475, B => N482, C => N474, Y => 
        ADD_27x27_fast_I213_Y_0);
    
    un2_resadd_ADD_27x27_fast_I16_P0N : OR2
      port map(A => ADDERinB(16), B => ADDERinA_16, Y => N374);
    
    \REG_RNO[16]\ : NOR2
      port map(A => clr_MAC_D, B => N_24, Y => \REG_4[16]\);
    
    un2_resadd_ADD_27x27_fast_I115_Y_0 : MIN3
      port map(A => ADDERinA_6, B => ADDERinB(6), C => N340, Y
         => ADD_27x27_fast_I115_Y_0);
    
    un2_resadd_ADD_27x27_fast_I47_Y : AO13
      port map(A => N367, B => ADDERinB(15), C => ADDERinA_15, Y
         => N425);
    
    \REG_RNO_0[0]\ : AX1E
      port map(A => ADDERinA_0, B => add_D_0, C => ADDERinB(0), Y
         => N_8);
    
    un2_resadd_ADD_27x27_fast_I114_Y : NOR2B
      port map(A => N446, B => N442, Y => N495);
    
    un2_resadd_ADD_27x27_fast_I251_Y_0 : AX1D
      port map(A => N415, B => ADD_27x27_fast_I210_Y_0_a2, C => 
        ADD_27x27_fast_I251_Y_0_0, Y => \un2_resadd[21]\);
    
    \REG_RNO[6]\ : NOR2
      port map(A => clr_MAC_D, B => N_14, Y => \REG_4[6]\);
    
    \REG_RNO[5]\ : NOR2
      port map(A => clr_MAC_D, B => N_13, Y => \REG_4[5]\);
    
    un2_resadd_ADD_27x27_fast_I56_Y : OA1
      port map(A => ADDERinA_11, B => ADDERinB(11), C => N356, Y
         => N434);
    
    \REG[2]\ : DFN1E0C0
      port map(D => \REG_4[2]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(2));
    
    un2_resadd_ADD_27x27_fast_I254_Y_0_0 : XOR2
      port map(A => ADDERinA_24, B => ADDERinB(24), Y => 
        ADD_27x27_fast_I254_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I10_P0N : OR2
      port map(A => ADDERinB(10), B => ADDERinA_10, Y => N356);
    
    \REG_RNO[23]\ : NOR2
      port map(A => clr_MAC_D, B => N_31, Y => \REG_4[23]\);
    
    un2_resadd_ADD_27x27_fast_I130_Y : NOR2
      port map(A => N471, B => N463, Y => N517);
    
    un2_resadd_ADD_27x27_fast_I209_Y_1 : OA1A
      port map(A => N474, B => N467, C => ADD_27x27_fast_I209_Y_0, 
        Y => ADD_27x27_fast_I209_Y_1);
    
    \REG[7]\ : DFN1E0C0
      port map(D => \REG_4[7]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(7));
    
    un2_resadd_ADD_27x27_fast_I211_Y_1 : AOI1B
      port map(A => N540, B => N525, C => ADD_27x27_fast_I211_Y_0, 
        Y => ADD_27x27_fast_I211_Y_1);
    
    un2_resadd_ADD_27x27_fast_I61_Y_0_o2 : AO1
      port map(A => N350, B => N346, C => N349, Y => N439);
    
    \REG_RNO[10]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_18, Y => \REG_4[10]\);
    
    \REG[4]\ : DFN1E0C0
      port map(D => \REG_4[4]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(4));
    
    \REG[10]\ : DFN1E0C0
      port map(D => \REG_4[10]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(10));
    
    un2_resadd_ADD_27x27_fast_I243_Y_0_0 : XOR2
      port map(A => ADDERinA_13, B => ADDERinB(13), Y => 
        ADD_27x27_fast_I243_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I208_Y_3 : AOI1B
      port map(A => N534, B => N519, C => ADD_27x27_fast_I208_Y_2, 
        Y => ADD_27x27_fast_I208_Y_3);
    
    un2_resadd_ADD_27x27_fast_I192_Y_0_a2 : OA1
      port map(A => I193_un1_Y, B => N540, C => N362, Y => 
        ADD_27x27_fast_I192_Y_0_a2);
    
    un2_resadd_ADD_27x27_fast_I190_Y : OR2
      port map(A => N534, B => I190_un1_Y, Y => N651);
    
    un2_resadd_ADD_27x27_fast_I18_P0N : OR2A
      port map(A => ADDERinA_i(18), B => ADDERinB(18), Y => N380);
    
    un2_resadd_ADD_27x27_fast_I207_un1_Y : OR3C
      port map(A => N533, B => N517, C => N548, Y => I207_un1_Y);
    
    un2_resadd_ADD_27x27_fast_I59_Y : MAJ3
      port map(A => ADDERinA_9, B => ADDERinB(9), C => N349, Y
         => N437);
    
    un2_resadd_ADD_27x27_fast_I251_Y_0_0 : XOR2
      port map(A => ADDERinA_21, B => ADDERinB(21), Y => 
        ADD_27x27_fast_I251_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I208_un1_Y : OR3C
      port map(A => N519, B => N535, C => N550, Y => I208_un1_Y);
    
    \REG_RNO[17]\ : NOR2
      port map(A => clr_MAC_D, B => N_25, Y => \REG_4[17]\);
    
    un1_clr_1 : NOR3
      port map(A => add_D_0, B => MACMUX2sel_D, C => clr_MAC_D_0, 
        Y => \un1_clr_1\);
    
    un2_resadd_ADD_27x27_fast_I98_Y : OR2B
      port map(A => N430, B => N426, Y => N479);
    
    un2_resadd_ADD_27x27_fast_I12_P0N : OR2
      port map(A => ADDERinB(12), B => ADDERinA_12, Y => N362);
    
    un2_resadd_ADD_27x27_fast_I117_Y : AO1
      port map(A => N449, B => N446, C => N445, Y => N498);
    
    un2_resadd_ADD_27x27_fast_I64_Y : OA1
      port map(A => ADDERinA_7, B => ADDERinB(7), C => N344, Y
         => N442);
    
    \REG[8]\ : DFN1E0C0
      port map(D => \REG_4[8]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(8));
    
    un2_resadd_ADD_27x27_fast_I240_Y_0 : AX1A
      port map(A => N544, B => I195_un1_Y_i, C => 
        ADD_27x27_fast_I240_Y_0_0, Y => \un2_resadd[10]\);
    
    un2_resadd_ADD_27x27_fast_I0_CO1 : OR2B
      port map(A => ADDERinB(0), B => ADDERinA_0, Y => N325);
    
    un2_resadd_ADD_27x27_fast_I34_Y : OA1
      port map(A => ADDERinA_21, B => ADDERinB(21), C => N392, Y
         => N412);
    
    un2_resadd_ADD_27x27_fast_I105_Y : AO1
      port map(A => N437, B => N434, C => N433, Y => N486);
    
    \REG_RNO_0[3]\ : MX2C
      port map(A => ADDERinB(3), B => \un2_resadd[3]\, S => 
        add_D_0, Y => N_11);
    
    un2_resadd_ADD_27x27_fast_I50_Y : OA1
      port map(A => ADDERinA_13, B => ADDERinB(13), C => N368, Y
         => N428);
    
    un2_resadd_ADD_27x27_fast_I239_Y_0 : AX1E
      port map(A => N_78_i, B => ADD_27x27_fast_I196_Y_0_0, C => 
        ADD_27x27_fast_I239_Y_0_0, Y => \un2_resadd[9]\);
    
    \REG[24]\ : DFN1E0C0
      port map(D => \REG_4[24]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(24));
    
    un2_resadd_ADD_27x27_fast_I3_P0N_i_o2 : OR2
      port map(A => ADDERinB(3), B => ADDERinA_3, Y => N_58);
    
    un2_resadd_ADD_27x27_fast_I15_P0N : OR2A
      port map(A => ADDERinA_15, B => ADDERinB(15), Y => N371);
    
    un2_resadd_ADD_27x27_fast_I249_Y_0 : AX1D
      port map(A => I212_un1_Y, B => ADD_27x27_fast_I212_Y_1, C
         => ADD_27x27_fast_I249_Y_0_0, Y => \un2_resadd[19]\);
    
    un2_resadd_ADD_27x27_fast_I189_Y : AOI1
      port map(A => N548, B => N533, C => N532, Y => N648_i);
    
    un2_resadd_ADD_27x27_fast_I4_G0N_i_o2 : NOR2B
      port map(A => ADDERinB(4), B => ADDERinA_4, Y => N_52_i_0);
    
    un2_resadd_ADD_27x27_fast_I250_Y_0_0 : XOR2
      port map(A => ADDERinA_20, B => ADDERinB(20), Y => 
        ADD_27x27_fast_I250_Y_0_0);
    
    \REG_RNO_0[12]\ : MX2C
      port map(A => ADDERinB(12), B => \un2_resadd[12]\, S => 
        add_D, Y => N_20);
    
    un2_resadd_ADD_27x27_fast_I44_Y : OA1
      port map(A => ADDERinA_17, B => ADDERinB(17), C => N374, Y
         => N422);
    
    un2_resadd_ADD_27x27_fast_I233_Y_0 : XOR3
      port map(A => ADDERinB(3), B => ADDERinA_3, C => N_48, Y
         => \un2_resadd[3]\);
    
    un2_resadd_ADD_27x27_fast_I194_un1_Y : OR2B
      port map(A => N_48, B => N543, Y => I194_un1_Y_i);
    
    un2_resadd_ADD_27x27_fast_I14_P0N : OR2A
      port map(A => ADDERinA_14, B => ADDERinB(14), Y => N368);
    
    un2_resadd_ADD_27x27_fast_I243_Y_0 : AX1A
      port map(A => ADD_27x27_fast_I192_Y_0_a2, B => N361, C => 
        ADD_27x27_fast_I243_Y_0_0, Y => \un2_resadd[13]\);
    
    un2_resadd_ADD_27x27_fast_I146_Y : NOR2
      port map(A => N487, B => N479, Y => N533);
    
    \REG_RNO_0[14]\ : MX2C
      port map(A => ADDERinB(14), B => \un2_resadd[14]\, S => 
        add_D_0, Y => N_22);
    
    \REG[16]\ : DFN1E0C0
      port map(D => \REG_4[16]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(16));
    
    un2_resadd_ADD_27x27_fast_I62_Y_i_o2 : OAI1
      port map(A => ADDERinA_7, B => ADDERinB(7), C => N350, Y
         => N_73);
    
    un2_resadd_ADD_27x27_fast_I210_Y_0_a2_1 : NOR2B
      port map(A => N386, B => N383, Y => N_105_1);
    
    un2_resadd_ADD_27x27_fast_I102_Y : OR2B
      port map(A => N434, B => N430, Y => N483);
    
    \REG_RNO_0[4]\ : MX2C
      port map(A => ADDERinB(4), B => \un2_resadd[4]\, S => 
        add_D_0, Y => N_12);
    
    un2_resadd_ADD_27x27_fast_I20_G0N : NOR2B
      port map(A => ADDERinB(20), B => ADDERinA_20, Y => N385);
    
    \REG_RNO_0[2]\ : MX2C
      port map(A => ADDERinB(2), B => \un2_resadd[2]\, S => add_D, 
        Y => N_10);
    
    un2_resadd_ADD_27x27_fast_I82_Y : OR2B
      port map(A => N414, B => N410, Y => N463);
    
    un2_resadd_ADD_27x27_fast_I234_Y_0 : XOR3
      port map(A => ADDERinB(4), B => ADDERinA_4, C => N502, Y
         => \un2_resadd[4]\);
    
    un2_resadd_ADD_27x27_fast_I250_Y_0 : AX1E
      port map(A => I211_un1_Y, B => ADD_27x27_fast_I211_Y_1, C
         => ADD_27x27_fast_I250_Y_0_0, Y => \un2_resadd[20]\);
    
    un2_resadd_ADD_27x27_fast_I252_Y_0_0 : XOR2
      port map(A => ADDERinA_22, B => ADDERinB(22), Y => 
        ADD_27x27_fast_I252_Y_0_0);
    
    un2_resadd_ADD_27x27_fast_I244_Y_0 : XOR3
      port map(A => ADDERinB(14), B => ADDERinA_14, C => N654_i, 
        Y => \un2_resadd[14]\);
    
    un2_resadd_ADD_27x27_fast_I69_Y_i_a2 : NOR2
      port map(A => N_59, B => N_52_i_0, Y => N_108);
    
    un2_resadd_ADD_27x27_fast_I18_G0N : NOR2A
      port map(A => ADDERinB(18), B => ADDERinA_i(18), Y => N379);
    
    un2_resadd_ADD_27x27_fast_I13_G0N : OR2B
      port map(A => ADDERinB(13), B => ADDERinA_13, Y => N364);
    
    \REG_RNO_0[5]\ : MX2C
      port map(A => ADDERinB(5), B => \un2_resadd[5]\, S => add_D, 
        Y => N_13);
    
    \REG[21]\ : DFN1E0C0
      port map(D => \REG_4[21]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1\, Q => ADDERout(21));
    
    un2_resadd_ADD_27x27_fast_I237_Y_0 : XOR3
      port map(A => ADDERinB(7), B => ADDERinA_7, C => N550, Y
         => \un2_resadd[7]\);
    
    \REG_RNO_0[22]\ : MX2C
      port map(A => ADDERinB(22), B => \un2_resadd[22]\, S => 
        add_D_0, Y => N_30);
    
    un2_resadd_ADD_27x27_fast_I107_Y : AO1B
      port map(A => N439, B => N436, C => ADD_27x27_fast_I107_Y_0, 
        Y => N488);
    
    un2_resadd_ADD_27x27_fast_I247_Y_0 : AX1A
      port map(A => N423, B => N_98_i, C => 
        ADD_27x27_fast_I247_Y_0_0, Y => \un2_resadd[17]\);
    
    \REG_RNO[0]\ : NOR2
      port map(A => clr_MAC_D_0, B => N_8, Y => \REG_4[0]\);
    
    \REG_RNO_0[15]\ : MX2C
      port map(A => ADDERinB(15), B => \un2_resadd[15]\, S => 
        add_D_0, Y => N_23);
    
    un2_resadd_ADD_27x27_fast_I148_Y : NOR2
      port map(A => N489, B => N481, Y => N535);
    
    \REG_RNO_0[24]\ : MX2C
      port map(A => ADDERinB(24), B => \un2_resadd[24]\, S => 
        add_D_0, Y => N_32);
    
    un2_resadd_ADD_27x27_fast_I253_Y_0 : AX1E
      port map(A => I208_un1_Y, B => ADD_27x27_fast_I208_Y_3, C
         => ADD_27x27_fast_I253_Y_0_0, Y => \un2_resadd[23]\);
    
    un2_resadd_ADD_27x27_fast_I213_un1_Y_0 : NOR3B
      port map(A => N499, B => N_47, C => N491, Y => 
        ADD_27x27_fast_I213_un1_Y_0);
    
    \REG[15]\ : DFN1E0C0
      port map(D => \REG_4[15]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \un1_clr_1_0\, Q => ADDERout(15));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_MUX2 is

    port( MULTout_D      : in    std_logic_vector(24 downto 7);
          ADDERout       : in    std_logic_vector(24 downto 7);
          sample_out_s   : out   std_logic_vector(17 downto 0);
          MACMUX2sel_D_D : in    std_logic
        );

end MAC_MUX2;

architecture DEF_ARCH of MAC_MUX2 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \RES[19]\ : MX2
      port map(A => ADDERout(19), B => MULTout_D(19), S => 
        MACMUX2sel_D_D, Y => sample_out_s(12));
    
    \RES[9]\ : MX2
      port map(A => ADDERout(9), B => MULTout_D(9), S => 
        MACMUX2sel_D_D, Y => sample_out_s(2));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \RES[12]\ : MX2
      port map(A => ADDERout(12), B => MULTout_D(12), S => 
        MACMUX2sel_D_D, Y => sample_out_s(5));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \RES[17]\ : MX2
      port map(A => ADDERout(17), B => MULTout_D(17), S => 
        MACMUX2sel_D_D, Y => sample_out_s(10));
    
    \RES[22]\ : MX2
      port map(A => ADDERout(22), B => MULTout_D(22), S => 
        MACMUX2sel_D_D, Y => sample_out_s(15));
    
    \RES[11]\ : MX2
      port map(A => ADDERout(11), B => MULTout_D(11), S => 
        MACMUX2sel_D_D, Y => sample_out_s(4));
    
    \RES[18]\ : MX2
      port map(A => ADDERout(18), B => MULTout_D(18), S => 
        MACMUX2sel_D_D, Y => sample_out_s(11));
    
    \RES[21]\ : MX2
      port map(A => ADDERout(21), B => MULTout_D(21), S => 
        MACMUX2sel_D_D, Y => sample_out_s(14));
    
    \RES[14]\ : MX2
      port map(A => ADDERout(14), B => MULTout_D(14), S => 
        MACMUX2sel_D_D, Y => sample_out_s(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \RES[24]\ : MX2
      port map(A => ADDERout(24), B => MULTout_D(24), S => 
        MACMUX2sel_D_D, Y => sample_out_s(17));
    
    \RES[10]\ : MX2
      port map(A => ADDERout(10), B => MULTout_D(10), S => 
        MACMUX2sel_D_D, Y => sample_out_s(3));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \RES[8]\ : MX2
      port map(A => ADDERout(8), B => MULTout_D(8), S => 
        MACMUX2sel_D_D, Y => sample_out_s(1));
    
    \RES[16]\ : MX2
      port map(A => ADDERout(16), B => MULTout_D(16), S => 
        MACMUX2sel_D_D, Y => sample_out_s(9));
    
    \RES[20]\ : MX2
      port map(A => ADDERout(20), B => MULTout_D(20), S => 
        MACMUX2sel_D_D, Y => sample_out_s(13));
    
    \RES[13]\ : MX2
      port map(A => ADDERout(13), B => MULTout_D(13), S => 
        MACMUX2sel_D_D, Y => sample_out_s(6));
    
    \RES[7]\ : MX2
      port map(A => ADDERout(7), B => MULTout_D(7), S => 
        MACMUX2sel_D_D, Y => sample_out_s(0));
    
    \RES[23]\ : MX2
      port map(A => ADDERout(23), B => MULTout_D(23), S => 
        MACMUX2sel_D_D, Y => sample_out_s(16));
    
    \RES[15]\ : MX2
      port map(A => ADDERout(15), B => MULTout_D(15), S => 
        MACMUX2sel_D_D, Y => sample_out_s(8));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC_REG_1_2 is

    port( MACMUXsel_D   : out   std_logic;
          MACMUXsel_D_0 : out   std_logic;
          N_4           : in    std_logic;
          HRESETn_c     : in    std_logic;
          HCLK_c        : in    std_logic;
          MACMUXsel_D_1 : out   std_logic
        );

end MAC_REG_1_2;

architecture DEF_ARCH of MAC_REG_1_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Q_1[0]\ : DFN1C0
      port map(D => N_4, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        MACMUXsel_D_1);
    
    \Q_0[0]\ : DFN1C0
      port map(D => N_4, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        MACMUXsel_D_0);
    
    \Q[0]\ : DFN1C0
      port map(D => N_4, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        MACMUXsel_D);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Multiplier is

    port( MULTout    : out   std_logic_vector(24 downto 0);
          alu_coef_s : in    std_logic_vector(8 downto 0);
          alu_sample : in    std_logic_vector(17 downto 0);
          mult       : in    std_logic;
          mult_0     : in    std_logic;
          HRESETn_c  : in    std_logic;
          HCLK_c     : in    std_logic
        );

end Multiplier;

architecture DEF_ARCH of Multiplier is 

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N399, ADD_22x22_fast_I80_un1_Y, N354, I120_un1_Y, 
        N407, N400, ADD_22x22_fast_I154_Y_0, 
        ADD_22x22_fast_I208_Y_0_0, N_253, N_250, 
        ADD_22x22_fast_I209_Y_0_2, N_252, 
        ADD_22x22_fast_I209_Y_0_0, N_254, \a17_b_i[7]\, 
        ADD_22x22_fast_I207_Y_0_0, N_249, N_244, 
        ADD_22x22_fast_I171_Y_2, I70_un1_Y, 
        ADD_22x22_fast_I171_Y_0, I110_un1_Y, N321, 
        ADD_22x22_fast_I206_Y_0_0, N_243, N_236, 
        ADD_22x22_fast_I170_Y_2, N395, N388, 
        ADD_22x22_fast_I170_Y_1, N346, N343, 
        ADD_22x22_fast_I170_Y_0, N324, ADD_22x22_fast_I205_Y_0_0, 
        madd_301, madd_527_0, N_235, ADD_22x22_fast_I172_Y_2, 
        I112_un1_Y, ADD_22x22_fast_I172_Y_0, I148_un1_Y, N350, 
        N347, ADD_22x22_fast_I200_Y_0_0, N_167, N_152, 
        ADD_22x22_fast_I203_Y_0_0, madd_262, madd_462_0, N_213, 
        ADD_22x22_fast_I173_Y_2, ADD_22x22_fast_I114_un1_Y, 
        ADD_22x22_fast_I173_Y_0, I173_un1_Y_i, 
        ADD_22x22_fast_I74_un1_Y, ADD_22x22_fast_I32_un1_Y, N318, 
        ADD_22x22_fast_I199_Y_0_0, N_134, N_149, N_136, 
        ADD_22x22_fast_I201_Y_0_0, N_150, N_165, N_183, 
        ADD_22x22_fast_I152_Y_0, N403, N396, 
        ADD_22x22_fast_I202_Y_0_0, N_182, madd_458_0_0, N_184, 
        ADD_22x22_fast_I198_Y_0_0, N_118, N_133, N_120, 
        ADD_22x22_fast_I172_un1_Y_0, N408, N416, N378, 
        ADD_22x22_fast_I153_un1_Y_0, N361, N398, N365, 
        ADD_22x22_fast_I155_Y_0, I82_un1_Y, N356, I155_un1_Y_i, 
        ADD_22x22_fast_I196_Y_0_0, N_86, N_101, N_88, 
        ADD_22x22_fast_I173_un1_Y_0, N410, N418, N_12, 
        ADD_22x22_fast_I152_un1_Y_0, I132_un1_Y_i, N411, N404, 
        ADD_22x22_fast_I197_Y_0_0, N_104, N_119, 
        ADD_22x22_fast_I157_un1_Y_0, N373, N421, N369, 
        ADD_22x22_fast_I155_un1_Y_0, I135_un1_Y_i, N417, 
        ADD_22x22_fast_I195_Y_0_0, N_72, N_87, 
        ADD_22x22_fast_I194_Y_0_0, N_69, madd_124_m6, N_56, 
        ADD_22x22_fast_I192_Y_0_0, N_28, N_39, N_30, N_180, 
        madd_458_14_0, N_195, madd_548_0_0, N_222, N_233, 
        ADD_22x22_fast_I190_Y_0_0, N_11_i, CO2, N_19, 
        madd_416_0_0, N_177_i, N_164, madd_268_0_0, N_113_i, 
        N_115, madd_522_0_tz_0, N_192, N_194, N_219, 
        madd_198_0_tz_0, N_61_i, N_63, N_50, madd_235_0_tz_0, 
        N_64_i, N_79, N_66, madd_24_0_0, N_7_i, N_9, 
        madd_120_0_0_1, N_32_i, N_43, N_34, madd_457_m5_0, N_185, 
        N_187, madd_39_0_0, N_15_i, N_13, madd_24_4_0, \a1_b[3]\, 
        \a0_b[4]\, madd_88_8_0, N_33_i, N_31, madd_268_8_0, 
        N_105_i, N_109, madd_115_0_0_1, \a0_b[8]\, \a2_b[6]\, 
        \a1_b[7]\, madd_493_6_0, \a_i10_b[8]\, madd_39_2_0, 
        \a5_b[0]\, \a3_b[2]\, madd_231_2_0, \a11_b[0]\, \a9_b[2]\, 
        madd_268_2_0, \a12_b[0]\, \a10_b[2]\, madd_523_4_0, 
        \a14_b[5]\, \a12_b[7]\, madd_458_2_0, madd_24_2_0, 
        \a2_b[2]\, \a4_b[0]\, madd_268_7_0, \a6_b[6]\, \a5_b[7]\, 
        madd_88_4_0, \a2_b[5]\, \a4_b[3]\, I157_un1_Y, I130_un1_Y, 
        ADD_22x22_fast_I171_un1_Y_0, madd_235_0_tz, N_99, N_174, 
        N_191, N402, I172_un1_Y, N392, ADD_22x22_fast_I115_Y_0, 
        I152_un1_Y, I154_un1_Y, N461, N_246_i, N_251, N_248, 
        \a16_b[7]\, \a_i15_b[8]\, \a17_b_i[6]\, N_240_i, N_247, 
        N_242, N_245, \a_i14_b[8]\, N_238, \a16_b[6]\, \a15_b[7]\, 
        \a17_b_i[5]\, N_241, N_239_i, N_234, N_237, \a16_b[5]\, 
        \a15_b[6]\, \a17_b_i[4]\, \a_i13_b[8]\, \a14_b[7]\, N_228, 
        N_230_i, N_232, N_224, N_231, N_229_i, N_220, N_227_i, 
        \a16_b[4]\, \a15_b[5]\, \a17_b_i[3]\, \a13_b[7]\, 
        \a14_b[6]\, \a_i12_b[8]\, N_218, N_216, N_225, N_223, 
        N_221, N_212, N_215, \a16_b[3]\, \a15_b[4]\, \a17_b_i[2]\, 
        N_217, \a13_b[6]\, N_204, \a_i11_b[8]\, N_202, N_208, 
        N_210, madd_457_m6, N_209_i, N_211, N_201, \a16_b[2]\, 
        \a15_b[3]\, \a17_b_i[1]\, N_203_i, \a12_b[6]\, \a14_b[4]\, 
        \a13_b[5]\, N_207, N_188_i, N_190, N_205, N_196, N_169_i, 
        \a15_b[1]\, \a16_b[0]\, \a14_b[2]\, N_171, \a11_b[5]\, 
        \a13_b[3]\, \a12_b[4]\, N_173, \a9_b[7]\, \a10_b[6]\, 
        \a_i8_b[8]\, N_175_i_0, N_156, N_154_i, N_158, N_163, 
        N_161_i, N_148, N_153_i, \a13_b[2]\, \a15_b[0]\, 
        \a14_b[1]\, N_155, \a10_b[5]\, \a12_b[3]\, \a11_b[4]\, 
        N_157, \a8_b[7]\, \a9_b[6]\, \a_i7_b[8]\, N_159_i, N_142, 
        N_138_i, N_140, N_146, N_144, N_147, N_145_i, N_132, 
        N_137_i, \a12_b[2]\, \a14_b[0]\, \a13_b[1]\, N_139, 
        \a9_b[5]\, \a11_b[3]\, \a10_b[4]\, N_141, \a_i6_b[8]\, 
        \a8_b[6]\, \a7_b[7]\, N_143_i, N_126, N_122_i, N_124, 
        N_130, N_128, N_131, N_129_i, N_116, N_121_i, \a11_b[2]\, 
        \a13_b[0]\, \a12_b[1]\, N_123, \a8_b[5]\, \a10_b[3]\, 
        \a9_b[4]\, N_125, \a6_b[7]\, \a7_b[6]\, \a_i5_b[8]\, 
        N_127_i, N_108, N_106_i, N_110, N_114, N_112, \a11_b[1]\, 
        N_107, \a7_b[5]\, \a9_b[3]\, \a8_b[4]\, \a_i4_b[8]\, 
        N_111_i, N_92, N_90_i, N_94, N_98, N_96, N_97, N_84, 
        N_89_i, \a10_b[1]\, N_91, \a6_b[5]\, \a8_b[3]\, \a7_b[4]\, 
        N_93, \a4_b[7]\, \a5_b[6]\, \a_i3_b[8]\, N_95_i, N_76, 
        N_74_i, N_78, N_82, N_80, N_85, N_83, N_81, N_68, N_73_i, 
        \a8_b[2]\, \a10_b[0]\, \a9_b[1]\, N_75, \a5_b[5]\, 
        \a7_b[3]\, \a6_b[4]\, N_77, \a4_b[6]\, \a_i2_b[8]\, 
        \a3_b[7]\, N_60, N_58_i, N_62, madd_119_m6, N_65_i, N_67, 
        N_57, \a7_b[2]\, \a9_b[0]\, \a8_b[1]\, N_59_i, \a5_b[4]\, 
        \a6_b[3]\, \a4_b[5]\, \a3_b[6]\, \a2_b[7]\, \a_i1_b[8]\, 
        N_44, \a_i0_b[8]\, N_46, N_48, N_45, \a3_b[5]\, \a5_b[3]\, 
        \a4_b[4]\, \a6_b[2]\, \a8_b[0]\, \a7_b[1]\, \a5_b[2]\, 
        \a7_b[0]\, \a6_b[1]\, \a3_b[4]\, N_37, N_24, N_25, N_14, 
        \a0_b[6]\, N_16, N_27, N_21_i, N_23, N_18, \a3_b[3]\, 
        \a2_b[4]\, \a1_b[5]\, N_17, N_8, \a4_b[1]\, \a0_b[5]\, 
        \a2_b[3]\, \a1_b[4]\, N_6, \a3_b[1]\, N_4, N_5, N_3, 
        \a0_b[3]\, N_2, \a3_b[0]\, \a2_b[1]\, \a1_b[2]\, N_1_i, 
        \a0_b[2]\, \a2_b[0]\, \a1_b[1]\, \a13_b[4]\, \a15_b[2]\, 
        \a14_b[3]\, N_189_i, \a10_b[7]\, \a12_b[5]\, \a11_b[6]\, 
        N_170, \a_i9_b[8]\, N_172, N_178, N_176, \RESMULT[24]\, 
        ADD_22x22_fast_I170_Y_3, \RESMULT[23]\, 
        ADD_22x22_fast_I171_Y_3, \RESMULT[22]\, \RESMULT[21]\, 
        I150_un1_Y, \RESMULT[20]\, \RESMULT[18]\, \RESMULT[17]\, 
        I122_un1_Y, \RESMULT[16]\, N449, I156_un1_Y_i, 
        \RESMULT[15]\, N451, \RESMULT[14]\, I158_un1_Y, N453, 
        \RESMULT[13]\, N455, I159_un1_Y_i, \RESMULT[12]\, 
        \RESMULT[10]\, \RESMULT[9]\, \RESMULT[8]\, N_53, N_55, 
        N419, \RESMULT[7]\, \RESMULT[6]\, N_29, \RESMULT[5]\, 
        \RESMULT[11]\, N413, I133_un1_Y_i, \RESMULT[19]\, N_214, 
        N544, \a17_b_i[0]\, N_186_1, N_206, I118_un1_Y, N397, 
        I153_un1_Y, N390, ADD_22x22_fast_I171_Y_3_tz, 
        ADD_22x22_fast_I170_Y_3_tz, N319, N313, N353, N349, 
        madd_61_2_0, \a6_b[0]\, \a5_b[1]\, N316, \a4_b[2]\, N_35, 
        \a0_b[7]\, \a1_b[6]\, N_22, madd_88_0_0, N_26, N_38, 
        N_40_i, N_51, N_36, N_179, N_162, N_160, madd_457_N_4, 
        madd_457tt_m3, madd_119_N_4, madd_119tt_m3, madd_124_N_4, 
        madd_124tt_m3, ADD_22x22_fast_I170_un1_Y_0, madd_462_0_tz, 
        madd_522_0, madd_487_0, madd_198_0, madd_477_0, 
        madd_477_0_tz, N412, madd_271, N_10, N_70, madd_112, 
        N_100, N_102, madd_133, N_166, madd_298, CO1, \a0_b[1]\, 
        \a1_b[0]\, \RESMULT[1]\, \RESMULT[2]\, \RESMULT[3]\, 
        \RESMULT[4]\, N273, N274, N276, N277, N279, N280, N288, 
        N289, N291, N292, N294, N295, N297, N298, N300, N301, 
        N303, N304, N306, N307, N352, N309, N312, N310, N357, 
        N362, N363, N364, N368, N285, N286, N372, N283, N376, 
        N377, N360, I90_un1_Y, N409, I101_un1_Y, N415, N345, N325, 
        N405, N282, N370, N374, N351, N358, N359, I92_un1_Y, N366, 
        N371, N375, I124_un1_Y, I134_un1_Y, madd_240, I126_un1_Y, 
        \RESMULT[0]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    RESMULT_madd_120_0 : XNOR3
      port map(A => N_38, B => madd_120_0_0_1, C => N_40_i, Y => 
        N_53);
    
    RESMULT_madd_452 : MIN3
      port map(A => N_189_i, B => N_176, C => N_178, Y => N_196);
    
    \RESMULT_a9_b[1]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(1), Y => 
        \a9_b[1]\);
    
    RESMULT_madd_65 : AO13
      port map(A => N_18, B => N_21_i, C => N_23, Y => N_28);
    
    RESMULT_madd_420 : AO18
      port map(A => N_164, B => N_179, C => N_177_i, Y => N_182);
    
    RESMULT_madd_606_ADD_22x22_fast_I3_P0N : OR2
      port map(A => N_55, B => N_53, Y => N283);
    
    RESMULT_madd_523_0 : XOR3
      port map(A => N_223, B => N_221, C => N_212, Y => N_225);
    
    \RESMULT_a4_b[2]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(2), Y => 
        \a4_b[2]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I124_un1_Y : NOR2B
      port map(A => N411, B => N404, Y => I124_un1_Y);
    
    RESMULT_madd_552 : MIN3
      port map(A => N_222, B => N_224, C => N_233, Y => N_236);
    
    \RESMULT_a9_b[4]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(4), Y => 
        \a9_b[4]\);
    
    RESMULT_madd_267 : MAJ3
      port map(A => N_111_i, B => N_96, C => N_98, Y => N_116);
    
    \RESMULT_a11_b[5]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(5), Y => 
        \a11_b[5]\);
    
    \RESMULT_a10_b[7]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(7), Y => 
        \a10_b[7]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I58_Y : AO1
      port map(A => N280, B => N276, C => N279, Y => N374);
    
    RESMULT_madd_606_ADD_22x22_fast_I55_Y : NOR2B
      port map(A => N286, B => N283, Y => N371);
    
    RESMULT_madd_606_ADD_22x22_fast_I99_Y : NOR2B
      port map(A => N377, B => N373, Y => N418);
    
    RESMULT_madd_606_ADD_22x22_fast_I156_un1_Y : OR3C
      port map(A => N404, B => N412, C => N419, Y => I156_un1_Y_i);
    
    RESMULT_madd_146 : MAJ3
      port map(A => \a_i0_b[8]\, B => N_44, C => N_46, Y => 
        N_64_i);
    
    RESMULT_madd_61_2_0 : XOR2
      port map(A => \a6_b[0]\, B => \a5_b[1]\, Y => madd_61_2_0);
    
    RESMULT_madd_378 : MAJ3
      port map(A => N_159_i, B => N_144, C => N_146, Y => N_164);
    
    RESMULT_madd_231_0 : XNOR3
      port map(A => N_99, B => N_97, C => N_84, Y => N_101);
    
    RESMULT_madd_606_ADD_22x22_fast_I173_Y_0 : NOR3A
      port map(A => ADD_22x22_fast_I74_un1_Y, B => 
        ADD_22x22_fast_I32_un1_Y, C => N318, Y => 
        ADD_22x22_fast_I173_Y_0);
    
    \RESMULT_a11_b[0]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(0), Y => 
        \a11_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I9_G0N : XA1A
      port map(A => N_134, B => N_149, C => N_136, Y => N300);
    
    \RESMULT_a13_b[7]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(7), Y => 
        \a13_b[7]\);
    
    RESMULT_madd_457_m5 : XOR3
      port map(A => N_174, B => madd_457_m5_0, C => N_191, Y => 
        madd_458_14_0);
    
    RESMULT_madd_43 : AO13
      port map(A => N_8, B => N_15_i, C => N_13, Y => N_18);
    
    RESMULT_madd_141 : MAJ3
      port map(A => \a3_b[6]\, B => \a2_b[7]\, C => \a_i1_b[8]\, 
        Y => N_62);
    
    \RESMULT_a7_b[7]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(7), Y => 
        \a7_b[7]\);
    
    RESMULT_madd_235 : AO1
      port map(A => madd_235_0_tz, B => N_97, C => madd_133, Y
         => N_102);
    
    RESMULT_madd_197 : NOR2A
      port map(A => N_83, B => N_68, Y => madd_112);
    
    RESMULT_madd_606_ADD_22x22_fast_I200_Y_0_0 : XOR2
      port map(A => N_167, B => N_152, Y => 
        ADD_22x22_fast_I200_Y_0_0);
    
    RESMULT_madd_38 : MIN3
      port map(A => \a2_b[3]\, B => \a0_b[5]\, C => \a1_b[4]\, Y
         => N_16);
    
    \REG[6]\ : DFN1E1C0
      port map(D => \RESMULT[6]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(6));
    
    RESMULT_madd_200 : NOR2A
      port map(A => N_85, B => N_70, Y => N_88);
    
    RESMULT_madd_104 : MAJ3
      port map(A => \a5_b[3]\, B => \a3_b[5]\, C => \a4_b[4]\, Y
         => N_46);
    
    \RESMULT_a14_b[7]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(7), Y => 
        \a14_b[7]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I31_Y : AO1C
      port map(A => N_243, B => N_236, C => N319, Y => N347);
    
    \RESMULT_a6_b[7]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(7), Y => 
        \a6_b[7]\);
    
    \RESMULT_a0_b[3]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(3), Y => 
        \a0_b[3]\);
    
    \RESMULT_a4_b[3]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(3), Y => 
        \a4_b[3]\);
    
    \RESMULT_a15_b[4]\ : NOR2B
      port map(A => alu_sample(15), B => alu_coef_s(4), Y => 
        \a15_b[4]\);
    
    RESMULT_madd_247 : MAJ3
      port map(A => \a9_b[3]\, B => \a7_b[5]\, C => \a8_b[4]\, Y
         => N_108);
    
    RESMULT_madd_606_ADD_22x22_fast_I172_un1_Y_0 : NOR3C
      port map(A => N408, B => N416, C => N378, Y => 
        ADD_22x22_fast_I172_un1_Y_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I122_un1_Y : OR2A
      port map(A => N409, B => N402, Y => I122_un1_Y);
    
    RESMULT_madd_523_8 : XOR3
      port map(A => N_217, B => N_215, C => N_206, Y => N_221);
    
    \RESMULT_a16_b[7]\ : OR2B
      port map(A => alu_sample(16), B => alu_coef_s(7), Y => 
        \a16_b[7]\);
    
    RESMULT_madd_457_m5_0 : XOR2
      port map(A => N_185, B => N_187, Y => madd_457_m5_0);
    
    RESMULT_madd_235_0_tz : OR2
      port map(A => madd_235_0_tz_0, B => N_99, Y => 
        madd_235_0_tz);
    
    RESMULT_madd_61_0 : XOR3
      port map(A => N_21_i, B => N_23, C => N_18, Y => N_27);
    
    \RESMULT_a9_b[0]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(0), Y => 
        \a9_b[0]\);
    
    \RESMULT_a6_b[1]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(1), Y => 
        \a6_b[1]\);
    
    \RESMULT_a13_b[0]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(0), Y => 
        \a13_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I73_Y : OR2A
      port map(A => N351, B => N347, Y => N392);
    
    RESMULT_madd_507 : MAJ3
      port map(A => \a14_b[5]\, B => \a12_b[7]\, C => \a13_b[6]\, 
        Y => N_218);
    
    RESMULT_madd_606_ADD_22x22_fast_I155_un1_Y : OR2A
      port map(A => ADD_22x22_fast_I155_un1_Y_0, B => N402, Y => 
        I155_un1_Y_i);
    
    RESMULT_madd_252 : MAJ3
      port map(A => \a6_b[6]\, B => \a5_b[7]\, C => \a_i4_b[8]\, 
        Y => N_110);
    
    RESMULT_madd_472 : MAJ3
      port map(A => \a14_b[4]\, B => \a12_b[6]\, C => \a13_b[5]\, 
        Y => N_204);
    
    RESMULT_madd_67 : NOR3B
      port map(A => N_17, B => N_25, C => N_10, Y => N_30);
    
    RESMULT_madd_95_0 : XNOR3
      port map(A => \a6_b[2]\, B => \a8_b[0]\, C => \a7_b[1]\, Y
         => N_43);
    
    \REG[18]\ : DFN1E1C0
      port map(D => \RESMULT[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(18));
    
    RESMULT_madd_568_4 : XOR3
      port map(A => \a_i13_b[8]\, B => \a14_b[7]\, C => N_228, Y
         => N_239_i);
    
    \RESMULT_a1_b[6]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(6), Y => 
        \a1_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I197_Y_0 : AX1A
      port map(A => N411, B => I132_un1_Y_i, C => 
        ADD_22x22_fast_I197_Y_0_0, Y => \RESMULT[12]\);
    
    RESMULT_madd_572 : AO18
      port map(A => N_234, B => N_241, C => N_239_i, Y => N_244);
    
    \RESMULT_a7_b[0]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(0), Y => 
        \a7_b[0]\);
    
    RESMULT_madd_88_4 : XOR2
      port map(A => madd_88_4_0, B => \a3_b[4]\, Y => N_33_i);
    
    RESMULT_madd_72 : MAJ3
      port map(A => \a7_b[0]\, B => \a5_b[2]\, C => \a6_b[1]\, Y
         => N_32_i);
    
    RESMULT_madd_230 : MAJ3
      port map(A => N_95_i, B => N_80, C => N_82, Y => N_100);
    
    RESMULT_madd_88_8 : XOR2
      port map(A => madd_88_8_0, B => N_24, Y => N_37);
    
    RESMULT_madd_606_ADD_22x22_fast_I80_un1_Y : NOR3C
      port map(A => N307, B => N310, C => N358, Y => 
        ADD_22x22_fast_I80_un1_Y);
    
    RESMULT_madd_458_0_0 : XNOR3
      port map(A => N_180, B => madd_458_14_0, C => N_195, Y => 
        madd_458_0_0);
    
    RESMULT_madd_66_0 : AX1
      port map(A => N_10, B => N_17, C => N_25, Y => N_29);
    
    RESMULT_madd_606_ADD_22x22_fast_I204_Y_0 : XOR3
      port map(A => N_225, B => N_214, C => N544, Y => 
        \RESMULT[19]\);
    
    RESMULT_madd_231_12 : XNOR3
      port map(A => N_82, B => N_95_i, C => N_80, Y => N_99);
    
    RESMULT_madd_194_4 : XNOR3
      port map(A => \a5_b[5]\, B => \a7_b[3]\, C => \a6_b[4]\, Y
         => N_75);
    
    RESMULT_madd_458_2 : XOR2
      port map(A => madd_458_2_0, B => \a17_b_i[0]\, Y => N_185);
    
    \RESMULT_a_i13_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(13), Y => 
        \a_i13_b[8]\);
    
    \REG[19]\ : DFN1E1C0
      port map(D => \RESMULT[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(19));
    
    \RESMULT_a6_b[0]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(0), Y => 
        \a6_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I34_Y : AO13
      port map(A => N312, B => N_225, C => N_214, Y => N350);
    
    RESMULT_madd_606_ADD_22x22_fast_I5_P0N : OR2
      port map(A => N_87, B => N_72, Y => N289);
    
    RESMULT_madd_606_ADD_22x22_fast_I197_Y_0_0 : XOR2
      port map(A => N_104, B => N_119, Y => 
        ADD_22x22_fast_I197_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I83_Y : OR2A
      port map(A => N361, B => N357, Y => N402);
    
    RESMULT_madd_537 : MAJ3
      port map(A => \a14_b[6]\, B => \a13_b[7]\, C => 
        \a_i12_b[8]\, Y => N_230_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I152_Y_0 : AO1
      port map(A => N403, B => N396, C => N395, Y => 
        ADD_22x22_fast_I152_Y_0);
    
    \RESMULT_a13_b[2]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(2), Y => 
        \a13_b[2]\);
    
    RESMULT_madd_416_4 : XNOR3
      port map(A => \a11_b[5]\, B => \a13_b[3]\, C => \a12_b[4]\, 
        Y => N_171);
    
    RESMULT_madd_606_ADD_22x22_fast_I42_Y : MAJ3
      port map(A => N_152, B => N_167, C => N300, Y => N358);
    
    RESMULT_madd_606_ADD_22x22_fast_I16_G0N : NOR2A
      port map(A => N_243, B => N_236, Y => N321);
    
    \RESMULT_a_i0_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(0), Y => 
        \a_i0_b[8]\);
    
    RESMULT_madd_437 : MAJ3
      port map(A => \a12_b[5]\, B => \a10_b[7]\, C => \a11_b[6]\, 
        Y => N_190);
    
    RESMULT_madd_606_ADD_22x22_fast_I100_Y : AO1
      port map(A => N378, B => N375, C => N374, Y => N419);
    
    RESMULT_madd_606_ADD_22x22_fast_I199_Y_0_0 : XNOR3
      port map(A => N_134, B => N_149, C => N_136, Y => 
        ADD_22x22_fast_I199_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I98_Y : AO1
      port map(A => N376, B => N373, C => N372, Y => N417);
    
    \RESMULT_a4_b[7]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(7), Y => 
        \a4_b[7]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I9_P0N : XO1A
      port map(A => N_134, B => N_149, C => N_136, Y => N301);
    
    RESMULT_madd_304 : MAJ3
      port map(A => N_127_i, B => N_112, C => N_114, Y => N_132);
    
    \RESMULT_a_i9_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(9), Y => 
        \a_i9_b[8]\);
    
    \REG[1]\ : DFN1E1C0
      port map(D => \RESMULT[1]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult_0, Q => MULTout(1));
    
    \RESMULT_a5_b[1]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(1), Y => 
        \a5_b[1]\);
    
    \RESMULT_a1_b[7]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(7), Y => 
        \a1_b[7]\);
    
    \RESMULT_a1_b[4]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(4), Y => 
        \a1_b[4]\);
    
    RESMULT_madd_476 : NOR2B
      port map(A => \a_i10_b[8]\, B => N_186_1, Y => madd_271);
    
    RESMULT_madd_39_2_0 : XOR2
      port map(A => \a5_b[0]\, B => \a3_b[2]\, Y => madd_39_2_0);
    
    RESMULT_madd_119_m6 : AO18
      port map(A => N_45, B => madd_115_0_0_1, C => madd_119_N_4, 
        Y => madd_119_m6);
    
    RESMULT_madd_606_ADD_22x22_fast_I133_un1_Y : OR3B
      port map(A => N373, B => N421, C => N369, Y => I133_un1_Y_i);
    
    RESMULT_madd_583_0 : XOR3
      port map(A => N_240_i, B => N_247, C => N_242, Y => N_249);
    
    RESMULT_madd_18 : MAJ3
      port map(A => \a4_b[0]\, B => \a2_b[2]\, C => \a3_b[1]\, Y
         => N_8);
    
    \RESMULT_a9_b[7]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(7), Y => 
        \a9_b[7]\);
    
    RESMULT_madd_492 : MAJ3
      port map(A => N_205, B => N_196, C => N_207, Y => N_212);
    
    \RESMULT_a0_b[5]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(5), Y => 
        \a0_b[5]\);
    
    \RESMULT_a2_b[4]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(4), Y => 
        \a2_b[4]\);
    
    RESMULT_madd_462_0 : NOR2B
      port map(A => madd_462_0_tz, B => N_195, Y => madd_462_0);
    
    RESMULT_madd_272 : AO13
      port map(A => N_100, B => N_113_i, C => N_115, Y => N_118);
    
    \RESMULT_a9_b[5]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(5), Y => 
        \a9_b[5]\);
    
    RESMULT_madd_225 : AO18
      port map(A => N_93, B => N_89_i, C => N_91, Y => N_98);
    
    RESMULT_madd_606_ADD_22x22_fast_I194_Y_0 : AX1A
      port map(A => N417, B => I135_un1_Y_i, C => 
        ADD_22x22_fast_I194_Y_0_0, Y => \RESMULT[9]\);
    
    RESMULT_madd_592 : MAJ3
      port map(A => \a_i15_b[8]\, B => \a16_b[7]\, C => 
        \a17_b_i[6]\, Y => N_252);
    
    RESMULT_madd_458_7 : XOR3
      port map(A => \a10_b[7]\, B => \a12_b[5]\, C => \a11_b[6]\, 
        Y => N_189_i);
    
    \RESMULT_a10_b[4]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(4), Y => 
        \a10_b[4]\);
    
    \RESMULT_a0_b[7]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(7), Y => 
        \a0_b[7]\);
    
    RESMULT_madd_588_0 : XNOR3
      port map(A => \a16_b[7]\, B => \a_i15_b[8]\, C => 
        \a17_b_i[6]\, Y => N_251);
    
    \RESMULT_a15_b[1]\ : OR2B
      port map(A => alu_sample(15), B => alu_coef_s(1), Y => 
        \a15_b[1]\);
    
    \RESMULT_a0_b[8]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(8), Y => 
        \a0_b[8]\);
    
    RESMULT_madd_24_4 : XNOR2
      port map(A => madd_24_4_0, B => N_4, Y => N_9);
    
    RESMULT_madd_606_ADD_22x22_fast_I198_Y_0 : AX1A
      port map(A => N455, B => I159_un1_Y_i, C => 
        ADD_22x22_fast_I198_Y_0_0, Y => \RESMULT[13]\);
    
    \REG[15]\ : DFN1E1C0
      port map(D => \RESMULT[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(15));
    
    RESMULT_madd_124_m2 : XOR2
      port map(A => N_37, B => N_35, Y => madd_88_0_0);
    
    \RESMULT_a_i5_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(5), Y => 
        \a_i5_b[8]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I134_Y : OR2
      port map(A => N415, B => I134_un1_Y, Y => N461);
    
    RESMULT_madd_606_ADD_22x22_fast_I8_P0N : XO1A
      port map(A => N_118, B => N_133, C => N_120, Y => N298);
    
    \REG[3]\ : DFN1E1C0
      port map(D => \RESMULT[3]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(3));
    
    RESMULT_madd_606_ADD_22x22_fast_I80_Y : OR2
      port map(A => ADD_22x22_fast_I80_un1_Y, B => N354, Y => 
        N399);
    
    RESMULT_madd_606_ADD_22x22_fast_I52_Y : MAJ3
      port map(A => N_72, B => N_87, C => N285, Y => N368);
    
    RESMULT_madd_606_ADD_22x22_fast_I27_Y : OA1
      port map(A => N_250, B => N_253, C => N325, Y => N343);
    
    \RESMULT_a_i12_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(12), Y => 
        \a_i12_b[8]\);
    
    RESMULT_madd_273_0 : XOR3
      port map(A => N_100, B => madd_268_0_0, C => N_102, Y => 
        N_119);
    
    \RESMULT_a10_b[6]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(6), Y => 
        \a10_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I71_Y : NOR2
      port map(A => N349, B => N345, Y => N390);
    
    RESMULT_madd_61_2 : XOR2
      port map(A => madd_61_2_0, B => \a4_b[2]\, Y => N_21_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I199_Y_0 : AX1D
      port map(A => I158_un1_Y, B => N453, C => 
        ADD_22x22_fast_I199_Y_0_0, Y => \RESMULT[14]\);
    
    \RESMULT_a6_b[5]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(5), Y => 
        \a6_b[5]\);
    
    RESMULT_madd_305_2 : XOR3
      port map(A => \a11_b[2]\, B => \a13_b[0]\, C => \a12_b[1]\, 
        Y => N_121_i);
    
    \RESMULT_a15_b[3]\ : OR2B
      port map(A => alu_sample(15), B => alu_coef_s(3), Y => 
        \a15_b[3]\);
    
    \RESMULT_a3_b[6]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(6), Y => 
        \a3_b[6]\);
    
    RESMULT_madd_342_2 : XOR3
      port map(A => \a12_b[2]\, B => \a14_b[0]\, C => \a13_b[1]\, 
        Y => N_137_i);
    
    \RESMULT_a5_b[6]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(6), Y => 
        \a5_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I172_Y_2 : NOR3C
      port map(A => I112_un1_Y, B => ADD_22x22_fast_I172_Y_0, C
         => I148_un1_Y, Y => ADD_22x22_fast_I172_Y_2);
    
    RESMULT_madd_331 : MAJ3
      port map(A => N_122_i, B => N_124, C => N_126, Y => N_144);
    
    RESMULT_madd_606_ADD_22x22_fast_I5_G0N : NOR2B
      port map(A => N_87, B => N_72, Y => N288);
    
    RESMULT_madd_606_ADD_22x22_fast_I171_Y_3 : OR3C
      port map(A => N398, B => N390, C => 
        ADD_22x22_fast_I171_Y_3_tz, Y => ADD_22x22_fast_I171_Y_3);
    
    RESMULT_madd_606_ADD_22x22_fast_I155_Y_0 : NOR3C
      port map(A => I82_un1_Y, B => N356, C => I155_un1_Y_i, Y
         => ADD_22x22_fast_I155_Y_0);
    
    RESMULT_madd_410 : AO18
      port map(A => N_173, B => N_169_i, C => N_171, Y => N_178);
    
    RESMULT_madd_220 : MAJ3
      port map(A => N_74_i, B => N_76, C => N_78, Y => N_96);
    
    RESMULT_madd_24_0 : XNOR2
      port map(A => madd_24_0_0, B => N_6, Y => N_11_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I6_G0N : XA1
      port map(A => N_86, B => N_101, C => N_88, Y => N291);
    
    RESMULT_madd_416_10 : XOR3
      port map(A => N_156, B => N_154_i, C => N_158, Y => 
        N_175_i_0);
    
    \RESMULT_a6_b[6]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(6), Y => 
        \a6_b[6]\);
    
    RESMULT_madd_363 : MAJ3
      port map(A => \a9_b[6]\, B => \a8_b[7]\, C => \a_i7_b[8]\, 
        Y => N_158);
    
    \RESMULT_a17_b_i[3]\ : NOR2A
      port map(A => alu_sample(17), B => alu_coef_s(3), Y => 
        \a17_b_i[3]\);
    
    \RESMULT_a8_b[2]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(2), Y => 
        \a8_b[2]\);
    
    RESMULT_madd_268_2 : XOR2
      port map(A => madd_268_2_0, B => \a11_b[1]\, Y => N_105_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I62_Y : AO1
      port map(A => N274, B => N_12, C => N273, Y => N378);
    
    \REG[10]\ : DFN1E1C0
      port map(D => \RESMULT[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(10));
    
    RESMULT_madd_606_ADD_22x22_fast_I135_un1_Y : OR2B
      port map(A => N418, B => N_12, Y => I135_un1_Y_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_Y_3_tz : OR2
      port map(A => N449, B => ADD_22x22_fast_I170_un1_Y_0, Y => 
        ADD_22x22_fast_I170_Y_3_tz);
    
    RESMULT_madd_194_0 : XNOR3
      port map(A => N_83, B => N_81, C => N_68, Y => N_85);
    
    RESMULT_madd_606_ADD_22x22_fast_I81_Y : OR3C
      port map(A => N307, B => N310, C => N359, Y => N400);
    
    \RESMULT_a11_b[6]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(6), Y => 
        \a11_b[6]\);
    
    \REG[12]\ : DFN1E1C0
      port map(D => \RESMULT[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(12));
    
    \RESMULT_a11_b[3]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(3), Y => 
        \a11_b[3]\);
    
    RESMULT_madd_55 : MAJ3
      port map(A => \a3_b[3]\, B => \a1_b[5]\, C => \a2_b[4]\, Y
         => N_24);
    
    \RESMULT_a_i4_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(4), Y => 
        \a_i4_b[8]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I6_P0N : XO1
      port map(A => N_86, B => N_101, C => N_88, Y => N292);
    
    RESMULT_madd_567 : AO13
      port map(A => N_232, B => N_230_i, C => N_237, Y => N_242);
    
    RESMULT_madd_421_0 : XOR3
      port map(A => N_179, B => madd_416_0_0, C => N_166, Y => 
        N_183);
    
    \RESMULT_a_i11_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(11), Y => 
        \a_i11_b[8]\);
    
    RESMULT_madd_342_12 : XNOR3
      port map(A => N_130, B => N_143_i, C => N_128, Y => N_147);
    
    RESMULT_madd_467 : MAJ3
      port map(A => \a15_b[3]\, B => \a16_b[2]\, C => 
        \a17_b_i[1]\, Y => N_202);
    
    RESMULT_madd_383 : AO13
      port map(A => N_148, B => N_161_i, C => N_163, Y => N_166);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_un1_Y_0 : NOR3C
      port map(A => N404, B => N412, C => N419, Y => 
        ADD_22x22_fast_I170_un1_Y_0);
    
    RESMULT_madd_379_0 : XOR3
      port map(A => N_163, B => N_161_i, C => N_148, Y => N_165);
    
    RESMULT_madd_606_ADD_22x22_fast_I46_Y : AO1
      port map(A => N298, B => N294, C => N297, Y => N362);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_Y_1 : AOI1B
      port map(A => N346, B => N343, C => ADD_22x22_fast_I170_Y_0, 
        Y => ADD_22x22_fast_I170_Y_1);
    
    RESMULT_madd_606_ADD_22x22_fast_I157_un1_Y_0 : NOR3B
      port map(A => N373, B => N421, C => N369, Y => 
        ADD_22x22_fast_I157_un1_Y_0);
    
    \REG[11]\ : DFN1E1C0
      port map(D => \RESMULT[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(11));
    
    RESMULT_madd_587 : AO18
      port map(A => N_242, B => N_247, C => N_240_i, Y => N_250);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \RESMULT_a7_b[3]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(3), Y => 
        \a7_b[3]\);
    
    \RESMULT_a8_b[6]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(6), Y => 
        \a8_b[6]\);
    
    \RESMULT_a3_b[3]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(3), Y => 
        \a3_b[3]\);
    
    RESMULT_madd_231_10 : XOR3
      port map(A => N_76, B => N_74_i, C => N_78, Y => N_95_i);
    
    RESMULT_madd_157_4 : XOR3
      port map(A => \a5_b[4]\, B => \a6_b[3]\, C => \a4_b[5]\, Y
         => N_59_i);
    
    RESMULT_madd_487 : MAJ3
      port map(A => N_203_i, B => N_192, C => N_194, Y => N_210);
    
    RESMULT_madd_157_9 : XNOR3
      port map(A => N_44, B => \a_i0_b[8]\, C => N_46, Y => N_63);
    
    RESMULT_madd_606_ADD_22x22_fast_I206_Y_0_0 : XNOR2
      port map(A => N_243, B => N_236, Y => 
        ADD_22x22_fast_I206_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I126_un1_Y : NOR3B
      port map(A => N361, B => N413, C => N365, Y => I126_un1_Y);
    
    RESMULT_madd_547 : AO13
      port map(A => N_220, B => N_229_i, C => N_231, Y => N_234);
    
    \RESMULT_a5_b[7]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(7), Y => 
        \a5_b[7]\);
    
    \REG[20]\ : DFN1E1C0
      port map(D => \RESMULT[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(20));
    
    RESMULT_madd_606_ADD_22x22_fast_I70_un1_Y : AO1D
      port map(A => N318, B => ADD_22x22_fast_I32_un1_Y, C => 
        N345, Y => I70_un1_Y);
    
    RESMULT_madd_60 : AO18
      port map(A => N_16, B => \a0_b[6]\, C => N_14, Y => N_26);
    
    \RESMULT_a10_b[0]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(0), Y => 
        \a10_b[0]\);
    
    \REG[22]\ : DFN1E1C0
      port map(D => \RESMULT[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult, Q => MULTout(22));
    
    RESMULT_madd_447 : MIN3
      port map(A => N_187, B => N_174, C => N_185, Y => N_194);
    
    RESMULT_madd_502 : MIN3
      port map(A => \a15_b[4]\, B => \a16_b[3]\, C => 
        \a17_b_i[2]\, Y => N_216);
    
    \RESMULT_a17_b_i[0]\ : OR2A
      port map(A => alu_sample(17), B => alu_coef_s(0), Y => 
        \a17_b_i[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I92_Y : OR2
      port map(A => N366, B => I92_un1_Y, Y => N411);
    
    RESMULT_madd_606_ADD_22x22_fast_I205_Y_0_0 : AX1B
      port map(A => madd_301, B => madd_527_0, C => N_235, Y => 
        ADD_22x22_fast_I205_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I84_Y : AO1
      port map(A => N362, B => N359, C => N358, Y => N403);
    
    RESMULT_madd_194_12 : XOR3
      port map(A => N_79, B => N_64_i, C => N_66, Y => N_83);
    
    \RESMULT_a15_b[0]\ : OR2B
      port map(A => alu_sample(15), B => alu_coef_s(0), Y => 
        \a15_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I190_Y_0 : XOR2
      port map(A => ADD_22x22_fast_I190_Y_0_0, B => N_12, Y => 
        \RESMULT[5]\);
    
    \RESMULT_a14_b[0]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(0), Y => 
        \a14_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I201_Y_0 : AX1A
      port map(A => N449, B => I156_un1_Y_i, C => 
        ADD_22x22_fast_I201_Y_0_0, Y => \RESMULT[16]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I155_un1_Y_0 : OA1A
      port map(A => I135_un1_Y_i, B => N417, C => N410, Y => 
        ADD_22x22_fast_I155_un1_Y_0);
    
    \REG[8]\ : DFN1E1C0
      port map(D => \RESMULT[8]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(8));
    
    RESMULT_madd_606_ADD_22x22_fast_I172_Y_0 : OA1C
      port map(A => N350, B => N347, C => N346, Y => 
        ADD_22x22_fast_I172_Y_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I11_G0N : NOR3B
      port map(A => N_165, B => N_183, C => N_150, Y => N306);
    
    \RESMULT_a16_b[3]\ : NOR2B
      port map(A => alu_sample(16), B => alu_coef_s(3), Y => 
        \a16_b[3]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I153_Y : NOR3
      port map(A => I118_un1_Y, B => N397, C => I153_un1_Y, Y => 
        N544);
    
    RESMULT_madd_606_ADD_22x22_fast_I191_Y_0 : XOR3
      port map(A => N_29, B => N_27, C => N378, Y => \RESMULT[6]\);
    
    \RESMULT_a5_b[3]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(3), Y => 
        \a5_b[3]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I38_Y : AO1
      port map(A => N310, B => N306, C => N309, Y => N354);
    
    RESMULT_madd_606_ADD_22x22_fast_I35_Y : NOR2B
      port map(A => N316, B => N313, Y => N351);
    
    RESMULT_madd_274 : XA1
      port map(A => N_100, B => madd_268_0_0, C => N_102, Y => 
        N_120);
    
    RESMULT_madd_606_ADD_22x22_fast_I56_Y : MAJ3
      port map(A => N_53, B => N_55, C => N279, Y => N372);
    
    RESMULT_madd_279 : MAJ3
      port map(A => \a13_b[0]\, B => \a11_b[2]\, C => \a12_b[1]\, 
        Y => N_122_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I10_G0N : NOR2B
      port map(A => N_167, B => N_152, Y => N303);
    
    \REG[21]\ : DFN1E1C0
      port map(D => \RESMULT[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult, Q => MULTout(21));
    
    RESMULT_madd_606_ADD_22x22_fast_I15_G0N : OA1
      port map(A => madd_301, B => madd_527_0, C => N_235, Y => 
        N318);
    
    RESMULT_madd_493_12 : XOR3
      port map(A => N_207, B => N_205, C => N_196, Y => N_211);
    
    RESMULT_madd_321 : MIN3
      port map(A => \a11_b[3]\, B => \a9_b[5]\, C => \a10_b[4]\, 
        Y => N_140);
    
    RESMULT_madd_342_7 : XNOR3
      port map(A => \a_i6_b[8]\, B => \a8_b[6]\, C => \a7_b[7]\, 
        Y => N_141);
    
    RESMULT_madd_432 : MAJ3
      port map(A => \a15_b[2]\, B => \a13_b[4]\, C => \a14_b[3]\, 
        Y => N_188_i);
    
    RESMULT_madd_268_7 : XNOR2
      port map(A => madd_268_7_0, B => \a_i4_b[8]\, Y => N_109);
    
    \REG[16]\ : DFN1E1C0
      port map(D => \RESMULT[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(16));
    
    RESMULT_madd_23 : MAJ3
      port map(A => \a1_b[3]\, B => N_4, C => \a0_b[4]\, Y => 
        N_10);
    
    \RESMULT_a14_b[4]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(4), Y => 
        \a14_b[4]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I82_un1_Y : OR2
      port map(A => N360, B => N357, Y => I82_un1_Y);
    
    RESMULT_madd_532 : MIN3
      port map(A => \a15_b[5]\, B => \a16_b[4]\, C => 
        \a17_b_i[3]\, Y => N_228);
    
    RESMULT_madd_24_2 : XOR2
      port map(A => madd_24_2_0, B => \a3_b[1]\, Y => N_7_i);
    
    \RESMULT_a16_b[4]\ : NOR2B
      port map(A => alu_sample(16), B => alu_coef_s(4), Y => 
        \a16_b[4]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I79_Y : NOR2
      port map(A => N357, B => N353, Y => N398);
    
    RESMULT_madd_606_ADD_22x22_fast_I17_P0N : OR2
      port map(A => N_249, B => N_244, Y => N325);
    
    RESMULT_madd_305_12 : XNOR3
      port map(A => N_114, B => N_127_i, C => N_112, Y => N_131);
    
    RESMULT_madd_543_4 : XOR3
      port map(A => \a13_b[7]\, B => \a14_b[6]\, C => 
        \a_i12_b[8]\, Y => N_229_i);
    
    \RESMULT_a14_b[3]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(3), Y => 
        \a14_b[3]\);
    
    \RESMULT_a_i6_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(6), Y => 
        \a_i6_b[8]\);
    
    \REG[4]\ : DFN1E1C0
      port map(D => \RESMULT[4]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(4));
    
    \REG[13]\ : DFN1E1C0
      port map(D => \RESMULT[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(13));
    
    RESMULT_madd_606_ADD_22x22_fast_I209_Y_0 : AX1E
      port map(A => ADD_22x22_fast_I170_Y_3, B => 
        ADD_22x22_fast_I170_Y_2, C => ADD_22x22_fast_I209_Y_0_2, 
        Y => \RESMULT[24]\);
    
    RESMULT_madd_336 : AO18
      port map(A => N_141, B => N_137_i, C => N_139, Y => N_146);
    
    RESMULT_madd_215 : MAJ3
      port map(A => \a5_b[6]\, B => \a4_b[7]\, C => \a_i3_b[8]\, 
        Y => N_94);
    
    RESMULT_madd_416_2 : XOR3
      port map(A => \a15_b[1]\, B => \a16_b[0]\, C => \a14_b[2]\, 
        Y => N_169_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I32_un1_Y : NOR3B
      port map(A => N_225, B => N319, C => N_214, Y => 
        ADD_22x22_fast_I32_un1_Y);
    
    RESMULT_madd_44_0 : XNOR2
      port map(A => N_17, B => N_10, Y => N_19);
    
    \RESMULT_a16_b[2]\ : OR2B
      port map(A => alu_sample(16), B => alu_coef_s(2), Y => 
        \a16_b[2]\);
    
    RESMULT_madd_341 : MAJ3
      port map(A => N_143_i, B => N_128, C => N_130, Y => N_148);
    
    \RESMULT_a17_b_i[5]\ : OR2A
      port map(A => alu_sample(17), B => alu_coef_s(5), Y => 
        \a17_b_i[5]\);
    
    RESMULT_madd_568_2 : XOR3
      port map(A => \a16_b[5]\, B => \a15_b[6]\, C => 
        \a17_b_i[4]\, Y => N_237);
    
    \RESMULT_a7_b[6]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(6), Y => 
        \a7_b[6]\);
    
    RESMULT_madd_305_7 : XNOR3
      port map(A => \a6_b[7]\, B => \a7_b[6]\, C => \a_i5_b[8]\, 
        Y => N_125);
    
    RESMULT_madd_606_ADD_22x22_fast_I0_P0N : AO1D
      port map(A => CO2, B => N_11_i, C => N_19, Y => N274);
    
    RESMULT_madd_606_ADD_22x22_fast_I2_G0N : XA1A
      port map(A => N_28, B => N_39, C => N_30, Y => N279);
    
    RESMULT_madd_606_ADD_22x22_fast_I89_Y : NOR3C
      port map(A => N289, B => N292, C => N363, Y => N408);
    
    RESMULT_madd_493_6_0 : AX1C
      port map(A => alu_coef_s(7), B => alu_sample(11), C => 
        \a_i10_b[8]\, Y => madd_493_6_0);
    
    RESMULT_madd_384_0 : XNOR2
      port map(A => N_165, B => N_150, Y => N_167);
    
    RESMULT_madd_305_0 : XOR3
      port map(A => N_131, B => N_129_i, C => N_116, Y => N_133);
    
    RESMULT_madd_294 : MAJ3
      port map(A => N_106_i, B => N_108, C => N_110, Y => N_128);
    
    RESMULT_madd_231_8 : XNOR3
      port map(A => N_91, B => N_89_i, C => N_93, Y => N_97);
    
    RESMULT_madd_268_2_0 : XOR2
      port map(A => \a12_b[0]\, B => \a10_b[2]\, Y => 
        madd_268_2_0);
    
    RESMULT_madd_299 : AO18
      port map(A => N_125, B => N_121_i, C => N_123, Y => N_130);
    
    RESMULT_madd_368 : AO18
      port map(A => N_142, B => N_138_i, C => N_140, Y => N_160);
    
    \RESMULT_a11_b[1]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(1), Y => 
        \a11_b[1]\);
    
    \REG[7]\ : DFN1E1C0
      port map(D => \RESMULT[7]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(7));
    
    RESMULT_madd_24_4_0 : XOR2
      port map(A => \a1_b[3]\, B => \a0_b[4]\, Y => madd_24_4_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I154_Y_0 : OR2
      port map(A => I120_un1_Y, B => N399, Y => 
        ADD_22x22_fast_I154_Y_0);
    
    \RESMULT_a5_b[2]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(2), Y => 
        \a5_b[2]\);
    
    RESMULT_madd_405 : MAJ3
      port map(A => N_154_i, B => N_156, C => N_158, Y => N_176);
    
    \RESMULT_a1_b[5]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(5), Y => 
        \a1_b[5]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I172_un1_Y : OR3A
      port map(A => ADD_22x22_fast_I172_un1_Y_0, B => N392, C => 
        N400, Y => I172_un1_Y);
    
    \REG[23]\ : DFN1E1C0
      port map(D => \RESMULT[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult, Q => MULTout(23));
    
    RESMULT_madd_606_ADD_22x22_fast_I10_P0N : OR2
      port map(A => N_167, B => N_152, Y => N304);
    
    RESMULT_madd_210 : MAJ3
      port map(A => \a8_b[3]\, B => \a6_b[5]\, C => \a7_b[4]\, Y
         => N_92);
    
    RESMULT_madd_114 : AO13
      port map(A => N_34, B => N_32_i, C => N_43, Y => N_50);
    
    \RESMULT_a12_b[0]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(0), Y => 
        \a12_b[0]\);
    
    \RESMULT_a_i15_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(15), Y => 
        \a_i15_b[8]\);
    
    \RESMULT_a7_b[5]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(5), Y => 
        \a7_b[5]\);
    
    RESMULT_madd_379_10 : XOR3
      port map(A => N_142, B => N_138_i, C => N_140, Y => N_159_i);
    
    RESMULT_madd_39_4 : XOR3
      port map(A => \a0_b[5]\, B => \a2_b[3]\, C => \a1_b[4]\, Y
         => N_15_i);
    
    \REG[0]\ : DFN1E1C0
      port map(D => \RESMULT[0]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult_0, Q => MULTout(0));
    
    RESMULT_madd_606_ADD_22x22_fast_I153_un1_Y_0 : NOR3B
      port map(A => N361, B => N398, C => N365, Y => 
        ADD_22x22_fast_I153_un1_Y_0);
    
    RESMULT_madd_458_9 : XNOR3
      port map(A => N_170, B => \a_i9_b[8]\, C => N_172, Y => 
        N_191);
    
    RESMULT_madd_606_ADD_22x22_fast_I101_Y : OR2
      port map(A => N376, B => I101_un1_Y, Y => N421);
    
    RESMULT_madd_157_11 : XNOR3
      port map(A => N_57, B => N_59_i, C => N_48, Y => N_65_i);
    
    \REG[5]\ : DFN1E1C0
      port map(D => \RESMULT[5]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(5));
    
    RESMULT_madd_606_ADD_22x22_fast_I114_un1_Y_0 : OR2
      port map(A => N353, B => N349, Y => ADD_22x22_fast_I115_Y_0);
    
    RESMULT_madd_125_0 : AX1
      port map(A => N_28, B => N_39, C => N_51, Y => N_55);
    
    \RESMULT_a8_b[1]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(1), Y => 
        \a8_b[1]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I96_Y : AO1
      port map(A => N374, B => N371, C => N370, Y => N415);
    
    RESMULT_madd_124tt_m3 : AO13
      port map(A => N_16, B => N_14, C => \a0_b[6]\, Y => 
        madd_124tt_m3);
    
    RESMULT_madd_493_8 : XOR3
      port map(A => N_188_i, B => N_201, C => N_190, Y => N_207);
    
    \RESMULT_a12_b[6]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(6), Y => 
        \a12_b[6]\);
    
    RESMULT_madd_348 : NOR2A
      port map(A => N_149, B => N_134, Y => N_152);
    
    RESMULT_madd_517 : MAJ3
      port map(A => N_215, B => N_206, C => N_217, Y => N_222);
    
    RESMULT_madd_606_ADD_22x22_fast_I207_Y_0_0 : XOR2
      port map(A => N_249, B => N_244, Y => 
        ADD_22x22_fast_I207_Y_0_0);
    
    \RESMULT_a12_b[7]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(7), Y => 
        \a12_b[7]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I173_Y_2 : NOR3C
      port map(A => ADD_22x22_fast_I114_un1_Y, B => 
        ADD_22x22_fast_I173_Y_0, C => I173_un1_Y_i, Y => 
        ADD_22x22_fast_I173_Y_2);
    
    \RESMULT_a12_b[3]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(3), Y => 
        \a12_b[3]\);
    
    RESMULT_madd_88_2 : XNOR3
      port map(A => \a5_b[2]\, B => \a7_b[0]\, C => \a6_b[1]\, Y
         => N_31);
    
    RESMULT_madd_523_7 : XNOR3
      port map(A => N_204, B => \a_i11_b[8]\, C => N_202, Y => 
        N_219);
    
    RESMULT_madd_422 : XO1
      port map(A => N_179, B => madd_416_0_0, C => N_166, Y => 
        N_184);
    
    RESMULT_madd_606_ADD_22x22_fast_I198_Y_0_0 : XNOR3
      port map(A => N_118, B => N_133, C => N_120, Y => 
        ADD_22x22_fast_I198_Y_0_0);
    
    RESMULT_madd_523_4_0 : XOR2
      port map(A => \a14_b[5]\, B => \a12_b[7]\, Y => 
        madd_523_4_0);
    
    \RESMULT_a4_b[5]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(5), Y => 
        \a4_b[5]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I47_Y : NOR2B
      port map(A => N298, B => N295, Y => N363);
    
    RESMULT_madd_606_ADD_22x22_fast_I110_un1_Y : OR2B
      port map(A => N397, B => N390, Y => I110_un1_Y);
    
    RESMULT_madd_548_0_0 : XOR2
      port map(A => N_222, B => N_233, Y => madd_548_0_0);
    
    RESMULT_madd_157_0 : XOR3
      port map(A => madd_119_m6, B => N_65_i, C => N_67, Y => 
        N_69);
    
    RESMULT_madd_606_ADD_22x22_fast_I78_Y : OAI1
      port map(A => N353, B => N356, C => N352, Y => N397);
    
    RESMULT_madd_522 : OR2
      port map(A => madd_522_0, B => madd_298, Y => N_224);
    
    RESMULT_madd_305_8 : XOR3
      port map(A => N_125, B => N_121_i, C => N_123, Y => N_129_i);
    
    RESMULT_madd_562 : MAJ3
      port map(A => \a14_b[7]\, B => N_228, C => \a_i13_b[8]\, Y
         => N_240_i);
    
    \REG[14]\ : DFN1E1C0
      port map(D => \RESMULT[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(14));
    
    \RESMULT_a2_b[6]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(6), Y => 
        \a2_b[6]\);
    
    \RESMULT_a0_b[1]\ : NOR2B
      port map(A => alu_sample(0), B => alu_coef_s(1), Y => 
        \a0_b[1]\);
    
    \RESMULT_a12_b[2]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(2), Y => 
        \a12_b[2]\);
    
    RESMULT_madd_157_7 : XOR3
      port map(A => \a3_b[6]\, B => \a2_b[7]\, C => \a_i1_b[8]\, 
        Y => N_61_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I11_P0N : AO1A
      port map(A => N_150, B => N_165, C => N_183, Y => N307);
    
    RESMULT_madd_1_605_SUM3_0 : XOR2
      port map(A => CO2, B => N_11_i, Y => \RESMULT[4]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I157_un1_Y : OR3B
      port map(A => N361, B => ADD_22x22_fast_I157_un1_Y_0, C => 
        N365, Y => I157_un1_Y);
    
    RESMULT_madd_178 : MAJ3
      port map(A => \a4_b[6]\, B => \a3_b[7]\, C => \a_i2_b[8]\, 
        Y => N_78);
    
    RESMULT_madd_326 : MIN3
      port map(A => \a8_b[6]\, B => \a7_b[7]\, C => \a_i6_b[8]\, 
        Y => N_142);
    
    RESMULT_madd_482 : AO18
      port map(A => N_190, B => N_201, C => N_188_i, Y => N_208);
    
    RESMULT_madd_606_ADD_22x22_fast_I171_Y_3_tz : OR2B
      port map(A => N451, B => ADD_22x22_fast_I171_un1_Y_0, Y => 
        ADD_22x22_fast_I171_Y_3_tz);
    
    RESMULT_madd_28 : AO18
      port map(A => N_6, B => N_9, C => N_7_i, Y => N_12);
    
    RESMULT_madd_606_ADD_22x22_fast_I150_un1_Y : OR3A
      port map(A => N455, B => ADD_22x22_fast_I115_Y_0, C => N402, 
        Y => I150_un1_Y);
    
    RESMULT_madd_582 : AO13
      port map(A => N_238, B => \a_i14_b[8]\, C => N_245, Y => 
        N_248);
    
    RESMULT_madd_543_2 : XNOR3
      port map(A => \a16_b[4]\, B => \a15_b[5]\, C => 
        \a17_b_i[3]\, Y => N_227_i);
    
    RESMULT_madd_194_8 : XNOR3
      port map(A => N_77, B => N_73_i, C => N_75, Y => N_81);
    
    \RESMULT_a17_b_i[1]\ : OR2A
      port map(A => alu_sample(17), B => alu_coef_s(1), Y => 
        \a17_b_i[1]\);
    
    \RESMULT_a0_b[4]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(4), Y => 
        \a0_b[4]\);
    
    RESMULT_madd_0_s : XOR3
      port map(A => \a0_b[2]\, B => \a2_b[0]\, C => \a1_b[1]\, Y
         => N_1_i);
    
    \RESMULT_a13_b[3]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(3), Y => 
        \a13_b[3]\);
    
    RESMULT_madd_442 : MAJ3
      port map(A => \a_i9_b[8]\, B => N_170, C => N_172, Y => 
        N_192);
    
    RESMULT_madd_606_ADD_22x22_fast_I90_un1_Y : NOR2A
      port map(A => N368, B => N365, Y => I90_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I88_Y : AO1
      port map(A => N366, B => N363, C => N362, Y => N407);
    
    RESMULT_madd_606_ADD_22x22_fast_I85_Y : NOR2B
      port map(A => N363, B => N359, Y => N404);
    
    RESMULT_madd_542 : MAJ3
      port map(A => N_227_i, B => N_216, C => N_218, Y => N_232);
    
    RESMULT_madd_522_0_tz_0 : OA1B
      port map(A => N_192, B => N_194, C => N_219, Y => 
        madd_522_0_tz_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I57_Y : NOR2B
      port map(A => N283, B => N280, Y => N373);
    
    \RESMULT_a4_b[6]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(6), Y => 
        \a4_b[6]\);
    
    \RESMULT_a0_b[2]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(2), Y => 
        \a0_b[2]\);
    
    RESMULT_madd_157_12 : XOR3
      port map(A => N_63, B => N_61_i, C => N_50, Y => N_67);
    
    \REG[24]\ : DFN1E1C0
      port map(D => \RESMULT[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult, Q => MULTout(24));
    
    RESMULT_madd_606_ADD_22x22_fast_I8_G0N : XA1A
      port map(A => N_118, B => N_133, C => N_120, Y => N297);
    
    RESMULT_madd_199_0 : XNOR2
      port map(A => N_85, B => N_70, Y => N_87);
    
    RESMULT_madd_50 : MAJ3
      port map(A => \a6_b[0]\, B => \a4_b[2]\, C => \a5_b[1]\, Y
         => N_22);
    
    RESMULT_madd_8 : MAJ3
      port map(A => \a3_b[0]\, B => \a1_b[2]\, C => \a2_b[1]\, Y
         => N_4);
    
    RESMULT_madd_477_0 : NOR3C
      port map(A => alu_coef_s(7), B => alu_sample(11), C => 
        madd_477_0_tz, Y => madd_477_0);
    
    RESMULT_madd_346 : AO13
      port map(A => N_132, B => N_145_i, C => N_147, Y => N_150);
    
    RESMULT_madd_262 : AO18
      port map(A => N_109, B => N_105_i, C => N_107, Y => N_114);
    
    RESMULT_madd_231_7 : XNOR3
      port map(A => \a4_b[7]\, B => \a5_b[6]\, C => \a_i3_b[8]\, 
        Y => N_93);
    
    RESMULT_madd_311 : NOR2A
      port map(A => N_133, B => N_118, Y => N_136);
    
    \RESMULT_a3_b[7]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(7), Y => 
        \a3_b[7]\);
    
    \RESMULT_a8_b[3]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(3), Y => 
        \a8_b[3]\);
    
    RESMULT_madd_173 : MAJ3
      port map(A => \a7_b[3]\, B => \a5_b[5]\, C => \a6_b[4]\, Y
         => N_76);
    
    \RESMULT_a14_b[6]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(6), Y => 
        \a14_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I4_P0N : XO1
      port map(A => N_69, B => madd_124_m6, C => N_56, Y => N286);
    
    RESMULT_madd_1_605_SUM2_0 : XOR2
      port map(A => CO1, B => N_5, Y => \RESMULT[3]\);
    
    RESMULT_madd_194_10 : XNOR3
      port map(A => N_60, B => N_58_i, C => N_62, Y => N_79);
    
    \RESMULT_a13_b[1]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(1), Y => 
        \a13_b[1]\);
    
    \RESMULT_a9_b[2]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(2), Y => 
        \a9_b[2]\);
    
    RESMULT_madd_198 : OR2
      port map(A => madd_198_0, B => madd_112, Y => N_86);
    
    RESMULT_madd_606_ADD_22x22_fast_I201_Y_0_0 : AX1
      port map(A => N_150, B => N_165, C => N_183, Y => 
        ADD_22x22_fast_I201_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I190_Y_0_0 : AX1B
      port map(A => N_11_i, B => CO2, C => N_19, Y => 
        ADD_22x22_fast_I190_Y_0_0);
    
    RESMULT_madd_156 : AO13
      port map(A => N_50, B => N_61_i, C => N_63, Y => N_68);
    
    RESMULT_madd_268_7_0 : XOR2
      port map(A => \a6_b[6]\, B => \a5_b[7]\, Y => madd_268_7_0);
    
    \RESMULT_a3_b[1]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(1), Y => 
        \a3_b[1]\);
    
    RESMULT_madd_268_10 : XOR3
      port map(A => N_92, B => N_90_i, C => N_94, Y => N_111_i);
    
    RESMULT_madd_342_4 : XNOR3
      port map(A => \a9_b[5]\, B => \a11_b[3]\, C => \a10_b[4]\, 
        Y => N_139);
    
    RESMULT_madd_606_ADD_22x22_fast_I7_P0N : OR2
      port map(A => N_119, B => N_104, Y => N295);
    
    RESMULT_madd_151 : AO13
      port map(A => N_48, B => N_59_i, C => N_57, Y => N_66);
    
    RESMULT_madd_606_ADD_22x22_fast_I209_Y_0_0 : AX1A
      port map(A => alu_sample(16), B => alu_coef_s(8), C => 
        \a17_b_i[7]\, Y => ADD_22x22_fast_I209_Y_0_0);
    
    \RESMULT_a12_b[5]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(5), Y => 
        \a12_b[5]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I206_Y_0 : AX1E
      port map(A => I150_un1_Y, B => ADD_22x22_fast_I173_Y_2, C
         => ADD_22x22_fast_I206_Y_0_0, Y => \RESMULT[21]\);
    
    \RESMULT_a17_b_i[4]\ : NOR2A
      port map(A => alu_sample(17), B => alu_coef_s(4), Y => 
        \a17_b_i[4]\);
    
    RESMULT_madd_234 : NOR2A
      port map(A => N_99, B => N_84, Y => madd_133);
    
    RESMULT_madd_99 : MAJ3
      port map(A => \a8_b[0]\, B => \a6_b[2]\, C => \a7_b[1]\, Y
         => N_44);
    
    RESMULT_madd_425 : NOR3C
      port map(A => alu_coef_s(1), B => alu_sample(16), C => 
        alu_sample(17), Y => madd_240);
    
    \RESMULT_a16_b[6]\ : OR2B
      port map(A => alu_sample(16), B => alu_coef_s(6), Y => 
        \a16_b[6]\);
    
    RESMULT_madd_242 : MAJ3
      port map(A => \a12_b[0]\, B => \a10_b[2]\, C => \a11_b[1]\, 
        Y => N_106_i);
    
    \RESMULT_a1_b[3]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(3), Y => 
        \a1_b[3]\);
    
    RESMULT_madd_521 : NOR2A
      port map(A => N_219, B => N_210, Y => madd_298);
    
    RESMULT_madd_606_ADD_22x22_fast_I13_G0N : OA1
      port map(A => madd_262, B => madd_462_0, C => N_213, Y => 
        N312);
    
    RESMULT_madd_568_6 : XOR3
      port map(A => N_237, B => N_230_i, C => N_232, Y => N_241);
    
    \RESMULT_a10_b[5]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(5), Y => 
        \a10_b[5]\);
    
    RESMULT_madd_124_m6 : MIN3
      port map(A => madd_120_0_0_1, B => madd_124_N_4, C => N_38, 
        Y => madd_124_m6);
    
    RESMULT_madd_606_ADD_22x22_fast_I205_Y_0 : AX1B
      port map(A => I152_un1_Y, B => ADD_22x22_fast_I152_Y_0, C
         => ADD_22x22_fast_I205_Y_0_0, Y => \RESMULT[20]\);
    
    RESMULT_madd_3 : MAJ3
      port map(A => \a2_b[0]\, B => \a0_b[2]\, C => \a1_b[1]\, Y
         => N_2);
    
    RESMULT_madd_379_4 : XNOR3
      port map(A => \a10_b[5]\, B => \a12_b[3]\, C => \a11_b[4]\, 
        Y => N_155);
    
    RESMULT_madd_257 : MAJ3
      port map(A => N_90_i, B => N_92, C => N_94, Y => N_112);
    
    RESMULT_madd_231_4 : XNOR3
      port map(A => \a6_b[5]\, B => \a8_b[3]\, C => \a7_b[4]\, Y
         => N_91);
    
    RESMULT_madd_115_2 : XNOR3
      port map(A => \a3_b[5]\, B => \a5_b[3]\, C => \a4_b[4]\, Y
         => N_45);
    
    RESMULT_madd_606_ADD_22x22_fast_I14_P0N : OR2A
      port map(A => N_214, B => N_225, Y => N316);
    
    RESMULT_madd_606_ADD_22x22_fast_I200_Y_0 : AX1E
      port map(A => I157_un1_Y, B => N451, C => 
        ADD_22x22_fast_I200_Y_0_0, Y => \RESMULT[15]\);
    
    \RESMULT_a2_b[1]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(1), Y => 
        \a2_b[1]\);
    
    RESMULT_madd_88_7 : XNOR3
      port map(A => \a0_b[7]\, B => \a1_b[6]\, C => N_22, Y => 
        N_35);
    
    RESMULT_madd_606_ADD_22x22_fast_I29_Y : AO1C
      port map(A => N_243, B => N_236, C => N325, Y => N345);
    
    RESMULT_madd_606_ADD_22x22_fast_I74_un1_Y : OR2
      port map(A => N352, B => N349, Y => 
        ADD_22x22_fast_I74_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I43_Y : NOR2B
      port map(A => N304, B => N301, Y => N359);
    
    RESMULT_madd_606_ADD_22x22_fast_I203_Y_0_0 : AX1B
      port map(A => madd_262, B => madd_462_0, C => N_213, Y => 
        ADD_22x22_fast_I203_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I173_un1_Y : OR3A
      port map(A => ADD_22x22_fast_I173_un1_Y_0, B => 
        ADD_22x22_fast_I115_Y_0, C => N402, Y => I173_un1_Y_i);
    
    RESMULT_madd_523_4 : XNOR2
      port map(A => madd_523_4_0, B => \a13_b[6]\, Y => N_217);
    
    RESMULT_madd_56_0 : XNOR3
      port map(A => N_14, B => \a0_b[6]\, C => N_16, Y => N_25);
    
    RESMULT_madd_606_ADD_22x22_fast_I13_P0N : OR3
      port map(A => madd_262, B => N_213, C => madd_462_0, Y => 
        N313);
    
    RESMULT_madd_193 : AO13
      port map(A => N_66, B => N_64_i, C => N_79, Y => N_84);
    
    RESMULT_madd_87 : AO13
      port map(A => N_24, B => N_33_i, C => N_31, Y => N_38);
    
    \RESMULT_a8_b[5]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(5), Y => 
        \a8_b[5]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I36_Y : AOI1
      port map(A => N313, B => N309, C => N312, Y => N352);
    
    RESMULT_madd_606_ADD_22x22_fast_I193_Y_0 : XOR3
      port map(A => N_53, B => N_55, C => N419, Y => \RESMULT[8]\);
    
    RESMULT_madd_1_605_CO2 : OR2B
      port map(A => CO1, B => N_5, Y => CO2);
    
    RESMULT_madd_606_ADD_22x22_fast_I97_Y : NOR2B
      port map(A => N375, B => N371, Y => N416);
    
    \RESMULT_a_i3_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(3), Y => 
        \a_i3_b[8]\);
    
    RESMULT_madd_124_m3 : MIN3
      port map(A => N_35, B => madd_124tt_m3, C => N_37, Y => 
        madd_124_N_4);
    
    \RESMULT_a16_b[5]\ : NOR2B
      port map(A => alu_sample(16), B => alu_coef_s(5), Y => 
        \a16_b[5]\);
    
    \RESMULT_a6_b[3]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(3), Y => 
        \a6_b[3]\);
    
    \RESMULT_a11_b[2]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(2), Y => 
        \a11_b[2]\);
    
    RESMULT_madd_462_0_tz : XO1A
      port map(A => N_180, B => madd_458_14_0, C => N_182, Y => 
        madd_462_0_tz);
    
    RESMULT_madd_493_2 : XNOR3
      port map(A => \a16_b[2]\, B => \a15_b[3]\, C => 
        \a17_b_i[1]\, Y => N_201);
    
    RESMULT_madd_606_ADD_22x22_fast_I130_un1_Y : NOR3A
      port map(A => N417, B => N369, C => N365, Y => I130_un1_Y);
    
    RESMULT_madd_268_0_0 : XOR2
      port map(A => N_113_i, B => N_115, Y => madd_268_0_0);
    
    \RESMULT_a3_b[5]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(5), Y => 
        \a3_b[5]\);
    
    \RESMULT_a2_b[5]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(5), Y => 
        \a2_b[5]\);
    
    \RESMULT_a16_b[0]\ : OR2B
      port map(A => alu_sample(16), B => alu_coef_s(0), Y => 
        \a16_b[0]\);
    
    RESMULT_madd_457tt_m3 : AO18
      port map(A => N_140, B => N_138_i, C => N_142, Y => 
        madd_457tt_m3);
    
    RESMULT_madd_194_2 : XOR3
      port map(A => \a8_b[2]\, B => \a10_b[0]\, C => \a9_b[1]\, Y
         => N_73_i);
    
    RESMULT_madd_457_m6 : MX2C
      port map(A => N_191, B => madd_457_N_4, S => madd_458_14_0, 
        Y => madd_457_m6);
    
    RESMULT_madd_305_10 : XOR3
      port map(A => N_108, B => N_106_i, C => N_110, Y => N_127_i);
    
    RESMULT_madd_9_0 : XOR3
      port map(A => N_3, B => \a0_b[3]\, C => N_2, Y => N_5);
    
    \REG[2]\ : DFN1E1C0
      port map(D => \RESMULT[2]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(2));
    
    RESMULT_madd_606_ADD_22x22_fast_I148_un1_Y : OR3A
      port map(A => N453, B => N392, C => N400, Y => I148_un1_Y);
    
    \REG[17]\ : DFN1E1C0
      port map(D => \RESMULT[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => mult_0, Q => MULTout(17));
    
    RESMULT_madd_606_ADD_22x22_fast_I53_Y : OR2B
      port map(A => N289, B => N286, Y => N369);
    
    RESMULT_madd_268_4 : XNOR3
      port map(A => \a7_b[5]\, B => \a9_b[3]\, C => \a8_b[4]\, Y
         => N_107);
    
    RESMULT_madd_231_2_0 : XOR2
      port map(A => \a11_b[0]\, B => \a9_b[2]\, Y => madd_231_2_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I195_Y_0_0 : XOR2
      port map(A => N_72, B => N_87, Y => 
        ADD_22x22_fast_I195_Y_0_0);
    
    RESMULT_madd_512 : MAJ3
      port map(A => \a_i11_b[8]\, B => N_202, C => N_204, Y => 
        N_220);
    
    RESMULT_madd_198_0_tz_0 : AO18
      port map(A => N_61_i, B => N_63, C => N_50, Y => 
        madd_198_0_tz_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I40_Y : AOI1
      port map(A => N307, B => N303, C => N306, Y => N356);
    
    RESMULT_madd_606_ADD_22x22_fast_I202_Y_0 : AX1E
      port map(A => I122_un1_Y, B => ADD_22x22_fast_I155_Y_0, C
         => ADD_22x22_fast_I202_Y_0_0, Y => \RESMULT[17]\);
    
    RESMULT_madd_120_0_0_1 : XNOR3
      port map(A => N_32_i, B => N_43, C => N_34, Y => 
        madd_120_0_0_1);
    
    RESMULT_madd_115_0 : XOR3
      port map(A => N_45, B => madd_115_0_0_1, C => N_36, Y => 
        N_51);
    
    RESMULT_madd_115_0_0_1 : XOR3
      port map(A => \a0_b[8]\, B => \a2_b[6]\, C => \a1_b[7]\, Y
         => madd_115_0_0_1);
    
    RESMULT_madd_493_4 : XOR3
      port map(A => \a12_b[6]\, B => \a14_b[4]\, C => \a13_b[5]\, 
        Y => N_203_i);
    
    RESMULT_madd_342_0 : XOR3
      port map(A => N_147, B => N_145_i, C => N_132, Y => N_149);
    
    RESMULT_madd_416_7 : XNOR3
      port map(A => \a9_b[7]\, B => \a10_b[6]\, C => \a_i8_b[8]\, 
        Y => N_173);
    
    RESMULT_madd_458_4 : XNOR3
      port map(A => \a13_b[4]\, B => \a15_b[2]\, C => \a14_b[3]\, 
        Y => N_187);
    
    \RESMULT_a9_b[6]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(6), Y => 
        \a9_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I1_P0N : OR2
      port map(A => N_29, B => N_27, Y => N277);
    
    \RESMULT_a14_b[2]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(2), Y => 
        \a14_b[2]\);
    
    RESMULT_madd_119_m3 : MIN3
      port map(A => \a0_b[7]\, B => madd_119tt_m3, C => \a1_b[6]\, 
        Y => madd_119_N_4);
    
    RESMULT_madd_523_10 : XNOR3
      port map(A => N_219, B => N_208, C => N_210, Y => N_223);
    
    RESMULT_madd_316 : MAJ3
      port map(A => \a14_b[0]\, B => \a12_b[2]\, C => \a13_b[1]\, 
        Y => N_138_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I192_Y_0_0 : XNOR3
      port map(A => N_28, B => N_39, C => N_30, Y => 
        ADD_22x22_fast_I192_Y_0_0);
    
    RESMULT_madd_88_8_0 : XOR2
      port map(A => N_33_i, B => N_31, Y => madd_88_8_0);
    
    \RESMULT_a14_b[1]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(1), Y => 
        \a14_b[1]\);
    
    \RESMULT_a15_b[6]\ : NOR2B
      port map(A => alu_sample(15), B => alu_coef_s(6), Y => 
        \a15_b[6]\);
    
    RESMULT_madd_342_8 : XOR3
      port map(A => N_141, B => N_137_i, C => N_139, Y => N_145_i);
    
    \RESMULT_a13_b[4]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(4), Y => 
        \a13_b[4]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I4_G0N : XA1
      port map(A => N_69, B => madd_124_m6, C => N_56, Y => N285);
    
    \RESMULT_a_i2_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(2), Y => 
        \a_i2_b[8]\);
    
    RESMULT_madd_39_2 : XNOR2
      port map(A => madd_39_2_0, B => \a4_b[1]\, Y => N_13);
    
    \RESMULT_a6_b[2]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(2), Y => 
        \a6_b[2]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I41_Y : OR2B
      port map(A => N307, B => N304, Y => N357);
    
    RESMULT_madd_606_ADD_22x22_fast_I50_Y : AO1
      port map(A => N292, B => N288, C => N291, Y => N366);
    
    RESMULT_madd_284 : MAJ3
      port map(A => \a10_b[3]\, B => \a8_b[5]\, C => \a9_b[4]\, Y
         => N_124);
    
    RESMULT_madd_606_ADD_22x22_fast_I152_un1_Y_0 : OA1A
      port map(A => I132_un1_Y_i, B => N411, C => N404, Y => 
        ADD_22x22_fast_I152_un1_Y_0);
    
    RESMULT_madd_289 : MAJ3
      port map(A => \a7_b[6]\, B => \a6_b[7]\, C => \a_i5_b[8]\, 
        Y => N_126);
    
    RESMULT_madd_606_ADD_22x22_fast_I209_Y_0_2 : XOR3
      port map(A => N_252, B => ADD_22x22_fast_I209_Y_0_0, C => 
        N_254, Y => ADD_22x22_fast_I209_Y_0_2);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_Y_0 : MIN3
      port map(A => N_250, B => N_253, C => N324, Y => 
        ADD_22x22_fast_I170_Y_0);
    
    \RESMULT_a3_b[0]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(0), Y => 
        \a3_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I171_un1_Y_0 : OR3B
      port map(A => N361, B => ADD_22x22_fast_I157_un1_Y_0, C => 
        N365, Y => ADD_22x22_fast_I171_un1_Y_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_Y_2 : AOI1B
      port map(A => N395, B => N388, C => ADD_22x22_fast_I170_Y_1, 
        Y => ADD_22x22_fast_I170_Y_2);
    
    \RESMULT_a7_b[1]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(1), Y => 
        \a7_b[1]\);
    
    RESMULT_madd_24_2_0 : XOR2
      port map(A => \a2_b[2]\, B => \a4_b[0]\, Y => madd_24_2_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I92_un1_Y : NOR3C
      port map(A => N289, B => N292, C => N370, Y => I92_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I114_un1_Y : AO1
      port map(A => N356, B => I82_un1_Y, C => 
        ADD_22x22_fast_I115_Y_0, Y => ADD_22x22_fast_I114_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I171_Y_0 : MIN3
      port map(A => N_244, B => N_249, C => N321, Y => 
        ADD_22x22_fast_I171_Y_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I124_Y : OR2
      port map(A => N403, B => I124_un1_Y, Y => N449);
    
    \RESMULT_a0_b[6]\ : OR2B
      port map(A => alu_sample(0), B => alu_coef_s(6), Y => 
        \a0_b[6]\);
    
    RESMULT_madd_523_2 : XOR3
      port map(A => \a16_b[3]\, B => \a15_b[4]\, C => 
        \a17_b_i[2]\, Y => N_215);
    
    RESMULT_madd_77 : MAJ3
      port map(A => \a4_b[3]\, B => \a2_b[5]\, C => \a3_b[4]\, Y
         => N_34);
    
    RESMULT_madd_606_ADD_22x22_fast_I2_P0N : XO1A
      port map(A => N_28, B => N_39, C => N_30, Y => N280);
    
    RESMULT_madd_157_2 : XNOR3
      port map(A => \a7_b[2]\, B => \a9_b[0]\, C => \a8_b[1]\, Y
         => N_57);
    
    RESMULT_madd_606_ADD_22x22_fast_I120_un1_Y : NOR2A
      port map(A => N407, B => N400, Y => I120_un1_Y);
    
    \RESMULT_a2_b[0]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(0), Y => 
        \a2_b[0]\);
    
    RESMULT_madd_379_7 : XNOR3
      port map(A => \a8_b[7]\, B => \a9_b[6]\, C => \a_i7_b[8]\, 
        Y => N_157);
    
    \RESMULT_a8_b[4]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(4), Y => 
        \a8_b[4]\);
    
    RESMULT_madd_461 : XA1A
      port map(A => N_180, B => madd_458_14_0, C => N_182, Y => 
        madd_262);
    
    \RESMULT_a2_b[3]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(3), Y => 
        \a2_b[3]\);
    
    \RESMULT_a17_b_i[6]\ : OR2A
      port map(A => alu_sample(17), B => alu_coef_s(6), Y => 
        \a17_b_i[6]\);
    
    \RESMULT_a12_b[1]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(1), Y => 
        \a12_b[1]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I76_Y : AO1
      port map(A => N354, B => N351, C => N350, Y => N395);
    
    RESMULT_madd_309 : AO13
      port map(A => N_116, B => N_129_i, C => N_131, Y => N_134);
    
    RESMULT_madd_1_605_SUM0_0 : XOR2
      port map(A => \a1_b[0]\, B => \a0_b[1]\, Y => \RESMULT[1]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I60_Y : MAJ3
      port map(A => N_27, B => N_29, C => N273, Y => N376);
    
    RESMULT_madd_606_ADD_22x22_fast_I154_un1_Y : NOR3B
      port map(A => N408, B => N461, C => N400, Y => I154_un1_Y);
    
    \RESMULT_a2_b[2]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(2), Y => 
        \a2_b[2]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I1_G0N : NOR2B
      port map(A => N_29, B => N_27, Y => N276);
    
    RESMULT_madd_415 : MAJ3
      port map(A => N_175_i_0, B => N_160, C => N_162, Y => N_180);
    
    RESMULT_madd_606_ADD_22x22_fast_I93_Y : NOR3C
      port map(A => N289, B => N292, C => N371, Y => N412);
    
    RESMULT_madd_543_0 : XOR3
      port map(A => N_231, B => N_229_i, C => N_220, Y => N_233);
    
    RESMULT_madd_119tt_m3 : MAJ3
      port map(A => \a6_b[0]\, B => \a4_b[2]\, C => \a5_b[1]\, Y
         => madd_119tt_m3);
    
    \RESMULT_a3_b[2]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(2), Y => 
        \a3_b[2]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I118_un1_Y : NOR2B
      port map(A => N405, B => N398, Y => I118_un1_Y);
    
    RESMULT_madd_493_11 : XOR3
      port map(A => N_192, B => N_203_i, C => N_194, Y => N_209_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I44_Y : AOI1
      port map(A => N301, B => N297, C => N300, Y => N360);
    
    RESMULT_madd_88_4_0 : XOR2
      port map(A => \a2_b[5]\, B => \a4_b[3]\, Y => madd_88_4_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I173_un1_Y_0 : NOR3C
      port map(A => N410, B => N418, C => N_12, Y => 
        ADD_22x22_fast_I173_un1_Y_0);
    
    \RESMULT_a9_b[3]\ : OR2B
      port map(A => alu_sample(9), B => alu_coef_s(3), Y => 
        \a9_b[3]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I171_Y_2 : NOR3C
      port map(A => I70_un1_Y, B => ADD_22x22_fast_I171_Y_0, C
         => I110_un1_Y, Y => ADD_22x22_fast_I171_Y_2);
    
    RESMULT_madd_606_ADD_22x22_fast_I112_un1_Y : AO1D
      port map(A => N354, B => ADD_22x22_fast_I80_un1_Y, C => 
        N392, Y => I112_un1_Y);
    
    RESMULT_madd_548_0 : XOR2
      port map(A => madd_548_0_0, B => N_224, Y => N_235);
    
    RESMULT_madd_606_ADD_22x22_fast_I196_Y_0_0 : XOR3
      port map(A => N_86, B => N_101, C => N_88, Y => 
        ADD_22x22_fast_I196_Y_0_0);
    
    \RESMULT_a4_b[4]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(4), Y => 
        \a4_b[4]\);
    
    \RESMULT_a15_b[7]\ : OR2B
      port map(A => alu_sample(15), B => alu_coef_s(7), Y => 
        \a15_b[7]\);
    
    RESMULT_madd_353 : MAJ3
      port map(A => \a15_b[0]\, B => \a13_b[2]\, C => \a14_b[1]\, 
        Y => N_154_i);
    
    \RESMULT_a_i10_b[8]\ : NOR2A
      port map(A => alu_coef_s(8), B => alu_sample(10), Y => 
        \a_i10_b[8]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I86_Y : AO1B
      port map(A => N364, B => N361, C => N360, Y => N405);
    
    RESMULT_madd_268_12 : XNOR3
      port map(A => N_98, B => N_111_i, C => N_96, Y => N_115);
    
    RESMULT_madd_1_605_CO1 : NOR3B
      port map(A => \a0_b[1]\, B => \a1_b[0]\, C => N_1_i, Y => 
        CO1);
    
    RESMULT_madd_4_0 : XNOR3
      port map(A => \a3_b[0]\, B => \a2_b[1]\, C => \a1_b[2]\, Y
         => N_3);
    
    \RESMULT_a17_b_i[2]\ : NOR2A
      port map(A => alu_sample(17), B => alu_coef_s(2), Y => 
        \a17_b_i[2]\);
    
    RESMULT_madd_379_12 : XNOR3
      port map(A => N_146, B => N_159_i, C => N_144, Y => N_163);
    
    RESMULT_madd_606_ADD_22x22_fast_I158_un1_Y : NOR3C
      port map(A => N408, B => N416, C => N378, Y => I158_un1_Y);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I37_Y : OR2B
      port map(A => N313, B => N310, Y => N353);
    
    RESMULT_madd_557 : MIN3
      port map(A => \a15_b[6]\, B => \a16_b[5]\, C => 
        \a17_b_i[4]\, Y => N_238);
    
    RESMULT_madd_458_13 : XNOR3
      port map(A => N_178, B => N_189_i, C => N_176, Y => N_195);
    
    RESMULT_madd_606_ADD_22x22_fast_I101_un1_Y : NOR2B
      port map(A => N377, B => N_12, Y => I101_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I159_un1_Y : OR3C
      port map(A => N410, B => N418, C => N_12, Y => I159_un1_Y_i);
    
    RESMULT_madd_457_m3 : MIN3
      port map(A => N_162, B => madd_457tt_m3, C => N_175_i_0, Y
         => madd_457_N_4);
    
    \RESMULT_a1_b[0]\ : NOR2B
      port map(A => alu_sample(1), B => alu_coef_s(0), Y => 
        \a1_b[0]\);
    
    RESMULT_madd_24_0_0 : XOR2
      port map(A => N_7_i, B => N_9, Y => madd_24_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I152_un1_Y : NOR2B
      port map(A => ADD_22x22_fast_I152_un1_Y_0, B => N396, Y => 
        I152_un1_Y);
    
    RESMULT_madd_606_ADD_22x22_fast_I17_G0N : NOR2B
      port map(A => N_249, B => N_244, Y => N324);
    
    RESMULT_madd_606_ADD_22x22_fast_I61_Y : NOR2B
      port map(A => N277, B => N274, Y => N377);
    
    RESMULT_madd_88_0 : XNOR2
      port map(A => madd_88_0_0, B => N_26, Y => N_39);
    
    RESMULT_madd_606_ADD_22x22_fast_I130_Y : OR2
      port map(A => N409, B => I130_un1_Y, Y => N455);
    
    RESMULT_madd_522_0 : OA1A
      port map(A => madd_522_0_tz_0, B => madd_487_0, C => N_208, 
        Y => madd_522_0);
    
    RESMULT_madd_487_0 : AOI1
      port map(A => N_194, B => N_192, C => N_203_i, Y => 
        madd_487_0);
    
    \RESMULT_a4_b[1]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(1), Y => 
        \a4_b[1]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I90_Y : OR2
      port map(A => N364, B => I90_un1_Y, Y => N409);
    
    \RESMULT_a13_b[6]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(6), Y => 
        \a13_b[6]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I54_Y : AO1
      port map(A => N286, B => N282, C => N285, Y => N370);
    
    \RESMULT_a2_b[7]\ : OR2B
      port map(A => alu_sample(2), B => alu_coef_s(7), Y => 
        \a2_b[7]\);
    
    RESMULT_madd_198_0 : OA1
      port map(A => N_83, B => madd_198_0_tz_0, C => N_81, Y => 
        madd_198_0);
    
    RESMULT_madd_168 : MAJ3
      port map(A => \a10_b[0]\, B => \a8_b[2]\, C => \a9_b[1]\, Y
         => N_74_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I196_Y_0 : AX1A
      port map(A => N413, B => I133_un1_Y_i, C => 
        ADD_22x22_fast_I196_Y_0_0, Y => \RESMULT[11]\);
    
    RESMULT_madd_109 : MAJ3
      port map(A => \a2_b[6]\, B => \a0_b[8]\, C => \a1_b[7]\, Y
         => N_48);
    
    \RESMULT_a10_b[2]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(2), Y => 
        \a10_b[2]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I126_Y : NOR2
      port map(A => N405, B => I126_un1_Y, Y => N451);
    
    \RESMULT_a17_b_i[7]\ : OR2A
      port map(A => alu_sample(17), B => alu_coef_s(7), Y => 
        \a17_b_i[7]\);
    
    RESMULT_madd_268_8_0 : XOR2
      port map(A => N_105_i, B => N_109, Y => madd_268_8_0);
    
    RESMULT_madd_573_0 : XNOR3
      port map(A => \a16_b[6]\, B => \a15_b[7]\, C => 
        \a17_b_i[5]\, Y => N_245);
    
    \RESMULT_a7_b[2]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(2), Y => 
        \a7_b[2]\);
    
    \RESMULT_a6_b[4]\ : OR2B
      port map(A => alu_sample(6), B => alu_coef_s(4), Y => 
        \a6_b[4]\);
    
    RESMULT_madd_92 : AO18
      port map(A => N_35, B => N_26, C => N_37, Y => N_40_i);
    
    RESMULT_madd_416_0_0 : XNOR2
      port map(A => N_177_i, B => N_164, Y => madd_416_0_0);
    
    RESMULT_madd_400 : MIN3
      port map(A => \a10_b[6]\, B => \a9_b[7]\, C => \a_i8_b[8]\, 
        Y => N_174);
    
    RESMULT_madd_390 : MAJ3
      port map(A => \a16_b[0]\, B => \a14_b[2]\, C => \a15_b[1]\, 
        Y => N_170);
    
    \RESMULT_a_i7_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(7), Y => 
        \a_i7_b[8]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I49_Y : OR2B
      port map(A => N295, B => N292, Y => N365);
    
    RESMULT_madd_606_ADD_22x22_fast_I12_G0N : XA1B
      port map(A => N_182, B => madd_458_0_0, C => N_184, Y => 
        N309);
    
    RESMULT_madd_458_2_0 : AX1E
      port map(A => alu_coef_s(1), B => alu_sample(16), C => 
        alu_sample(17), Y => madd_458_2_0);
    
    RESMULT_madd_568_0 : XOR3
      port map(A => N_241, B => N_239_i, C => N_234, Y => N_243);
    
    RESMULT_madd_527_0 : OA1
      port map(A => N_212, B => N_223, C => N_221, Y => 
        madd_527_0);
    
    RESMULT_madd_526 : NOR2B
      port map(A => N_223, B => N_212, Y => madd_301);
    
    RESMULT_madd_427_1 : OR2A
      port map(A => \a17_b_i[0]\, B => madd_240, Y => N_186_1);
    
    RESMULT_madd_188 : AO18
      port map(A => N_77, B => N_73_i, C => N_75, Y => N_82);
    
    \RESMULT_a8_b[7]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(7), Y => 
        \a8_b[7]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I15_P0N : OR3
      port map(A => N_235, B => madd_301, C => madd_527_0, Y => 
        N319);
    
    RESMULT_madd_543_6 : XNOR3
      port map(A => N_218, B => N_227_i, C => N_216, Y => N_231);
    
    RESMULT_madd_136 : MAJ3
      port map(A => \a6_b[3]\, B => \a4_b[5]\, C => \a5_b[4]\, Y
         => N_60);
    
    \RESMULT_a3_b[4]\ : OR2B
      port map(A => alu_sample(3), B => alu_coef_s(4), Y => 
        \a3_b[4]\);
    
    RESMULT_madd_373 : AO18
      port map(A => N_157, B => N_153_i, C => N_155, Y => N_162);
    
    RESMULT_madd_578_0 : XOR3
      port map(A => N_245, B => \a_i14_b[8]\, C => N_238, Y => 
        N_247);
    
    \RESMULT_a5_b[5]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(5), Y => 
        \a5_b[5]\);
    
    \RESMULT_a15_b[5]\ : NOR2B
      port map(A => alu_sample(15), B => alu_coef_s(5), Y => 
        \a15_b[5]\);
    
    RESMULT_madd_231_2 : XOR2
      port map(A => madd_231_2_0, B => \a10_b[1]\, Y => N_89_i);
    
    \RESMULT_a5_b[0]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(0), Y => 
        \a5_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I91_Y : NOR2
      port map(A => N369, B => N365, Y => N410);
    
    RESMULT_madd_477_0_tz : OR2
      port map(A => \a_i10_b[8]\, B => N_186_1, Y => 
        madd_477_0_tz);
    
    RESMULT_madd_131 : MAJ3
      port map(A => \a9_b[0]\, B => \a7_b[2]\, C => \a8_b[1]\, Y
         => N_58_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I128_Y : AO1
      port map(A => N415, B => N408, C => N407, Y => N453);
    
    RESMULT_madd_577 : MAJ3
      port map(A => \a15_b[7]\, B => \a16_b[6]\, C => 
        \a17_b_i[5]\, Y => N_246_i);
    
    RESMULT_madd_305_4 : XNOR3
      port map(A => \a8_b[5]\, B => \a10_b[3]\, C => \a9_b[4]\, Y
         => N_123);
    
    RESMULT_madd_61_4 : XNOR3
      port map(A => \a3_b[3]\, B => \a2_b[4]\, C => \a1_b[5]\, Y
         => N_23);
    
    RESMULT_madd_477 : OR2
      port map(A => madd_477_0, B => madd_271, Y => N_206);
    
    RESMULT_madd_416_12 : XNOR3
      port map(A => N_162, B => N_175_i_0, C => N_160, Y => N_179);
    
    RESMULT_madd_606_ADD_22x22_fast_I192_Y_0 : XOR2
      port map(A => ADD_22x22_fast_I192_Y_0_0, B => N421, Y => 
        \RESMULT[7]\);
    
    RESMULT_madd_194_7 : XNOR3
      port map(A => \a4_b[6]\, B => \a_i2_b[8]\, C => \a3_b[7]\, 
        Y => N_77);
    
    RESMULT_madd_163 : NOR2B
      port map(A => madd_124_m6, B => N_69, Y => N_72);
    
    \RESMULT_a13_b[5]\ : OR2B
      port map(A => alu_sample(13), B => alu_coef_s(5), Y => 
        \a13_b[5]\);
    
    \RESMULT_a1_b[1]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(1), Y => 
        \a1_b[1]\);
    
    RESMULT_madd_237 : NOR2B
      port map(A => N_101, B => N_86, Y => N_104);
    
    RESMULT_madd_593_0 : XOR3
      port map(A => N_246_i, B => N_251, C => N_248, Y => N_253);
    
    RESMULT_madd_379_2 : XOR3
      port map(A => \a13_b[2]\, B => \a15_b[0]\, C => \a14_b[1]\, 
        Y => N_153_i);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I3_G0N : NOR2B
      port map(A => N_55, B => N_53, Y => N282);
    
    RESMULT_madd_606_ADD_22x22_fast_I134_un1_Y : NOR2B
      port map(A => N416, B => N378, Y => I134_un1_Y);
    
    RESMULT_madd_493_0 : XOR3
      port map(A => madd_457_m6, B => N_209_i, C => N_211, Y => 
        N_213);
    
    RESMULT_madd_33 : MIN3
      port map(A => \a5_b[0]\, B => \a3_b[2]\, C => \a4_b[1]\, Y
         => N_14);
    
    RESMULT_madd_606_ADD_22x22_fast_I59_Y : NOR2B
      port map(A => N280, B => N277, Y => N375);
    
    \RESMULT_a8_b[0]\ : OR2B
      port map(A => alu_sample(8), B => alu_coef_s(0), Y => 
        \a8_b[0]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I202_Y_0_0 : XNOR3
      port map(A => N_182, B => madd_458_0_0, C => N_184, Y => 
        ADD_22x22_fast_I202_Y_0_0);
    
    RESMULT_madd_183 : MAJ3
      port map(A => N_58_i, B => N_60, C => N_62, Y => N_80);
    
    RESMULT_madd_606_ADD_22x22_fast_I0_G0N : NOR3A
      port map(A => N_19, B => N_11_i, C => CO2, Y => N273);
    
    \RESMULT_a11_b[4]\ : OR2B
      port map(A => alu_sample(11), B => alu_coef_s(4), Y => 
        \a11_b[4]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I170_Y_3 : OR3C
      port map(A => N396, B => N388, C => 
        ADD_22x22_fast_I170_Y_3_tz, Y => ADD_22x22_fast_I170_Y_3);
    
    RESMULT_madd_606_ADD_22x22_fast_I94_Y : AO1A
      port map(A => N369, B => N372, C => N368, Y => N413);
    
    RESMULT_madd_606_ADD_22x22_fast_I77_Y : NOR3C
      port map(A => N307, B => N310, C => N351, Y => N396);
    
    \RESMULT_a0_b[0]\ : NOR2B
      port map(A => alu_sample(0), B => alu_coef_s(0), Y => 
        \RESMULT[0]\);
    
    RESMULT_madd_39_0 : XOR2
      port map(A => madd_39_0_0, B => N_8, Y => N_17);
    
    RESMULT_madd_606_ADD_22x22_fast_I33_Y : OR2B
      port map(A => N319, B => N316, Y => N349);
    
    RESMULT_madd_606_ADD_22x22_fast_I208_Y_0 : AX1E
      port map(A => ADD_22x22_fast_I171_Y_3, B => 
        ADD_22x22_fast_I171_Y_2, C => ADD_22x22_fast_I208_Y_0_0, 
        Y => \RESMULT[23]\);
    
    \RESMULT_a_i1_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(1), Y => 
        \a_i1_b[8]\);
    
    RESMULT_madd_39_0_0 : XOR2
      port map(A => N_15_i, B => N_13, Y => madd_39_0_0);
    
    RESMULT_madd_342_10 : XOR3
      port map(A => N_126, B => N_122_i, C => N_124, Y => N_143_i);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    RESMULT_madd_597 : AO13
      port map(A => N_248, B => N_246_i, C => N_251, Y => N_254);
    
    \RESMULT_a7_b[4]\ : OR2B
      port map(A => alu_sample(7), B => alu_coef_s(4), Y => 
        \a7_b[4]\);
    
    RESMULT_madd_358 : MAJ3
      port map(A => \a12_b[3]\, B => \a10_b[5]\, C => \a11_b[4]\, 
        Y => N_156);
    
    RESMULT_madd_235_0_tz_0 : AO18
      port map(A => N_64_i, B => N_79, C => N_66, Y => 
        madd_235_0_tz_0);
    
    \RESMULT_a10_b[1]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(1), Y => 
        \a10_b[1]\);
    
    RESMULT_madd_497 : AO13
      port map(A => madd_457_m6, B => N_209_i, C => N_211, Y => 
        N_214);
    
    RESMULT_madd_395 : MAJ3
      port map(A => \a13_b[3]\, B => \a11_b[5]\, C => \a12_b[4]\, 
        Y => N_172);
    
    \RESMULT_a10_b[3]\ : OR2B
      port map(A => alu_sample(10), B => alu_coef_s(3), Y => 
        \a10_b[3]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I208_Y_0_0 : XOR2
      port map(A => N_253, B => N_250, Y => 
        ADD_22x22_fast_I208_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I69_Y : NOR2A
      port map(A => N343, B => N347, Y => N388);
    
    RESMULT_madd_606_ADD_22x22_fast_I132_un1_Y : OR2B
      port map(A => N419, B => N412, Y => I132_un1_Y_i);
    
    RESMULT_madd_268_8 : XOR2
      port map(A => madd_268_8_0, B => N_107, Y => N_113_i);
    
    RESMULT_madd_1_605_SUM1_0 : AX1E
      port map(A => \a0_b[1]\, B => \a1_b[0]\, C => N_1_i, Y => 
        \RESMULT[2]\);
    
    \REG[9]\ : DFN1E1C0
      port map(D => \RESMULT[9]\, CLK => HCLK_c, CLR => HRESETn_c, 
        E => mult, Q => MULTout(9));
    
    RESMULT_madd_606_ADD_22x22_fast_I203_Y_0 : AX1B
      port map(A => I154_un1_Y, B => ADD_22x22_fast_I154_Y_0, C
         => ADD_22x22_fast_I203_Y_0_0, Y => \RESMULT[18]\);
    
    \RESMULT_a15_b[2]\ : OR2B
      port map(A => alu_sample(15), B => alu_coef_s(2), Y => 
        \a15_b[2]\);
    
    RESMULT_madd_379_8 : XOR3
      port map(A => N_155, B => N_153_i, C => N_157, Y => N_161_i);
    
    RESMULT_madd_82 : MAJ3
      port map(A => \a1_b[6]\, B => N_22, C => \a0_b[7]\, Y => 
        N_36);
    
    RESMULT_madd_606_ADD_22x22_fast_I48_Y : MAJ3
      port map(A => N_104, B => N_119, C => N291, Y => N364);
    
    RESMULT_madd_606_ADD_22x22_fast_I45_Y : NOR2B
      port map(A => N301, B => N298, Y => N361);
    
    \RESMULT_a5_b[4]\ : OR2B
      port map(A => alu_sample(5), B => alu_coef_s(4), Y => 
        \a5_b[4]\);
    
    RESMULT_madd_416_8 : XOR3
      port map(A => N_171, B => N_169_i, C => N_173, Y => N_177_i);
    
    RESMULT_madd_606_ADD_22x22_fast_I12_P0N : XAI1A
      port map(A => N_182, B => madd_458_0_0, C => N_184, Y => 
        N310);
    
    RESMULT_madd_606_ADD_22x22_fast_I195_Y_0 : XOR2
      port map(A => ADD_22x22_fast_I195_Y_0_0, B => N461, Y => 
        \RESMULT[10]\);
    
    \RESMULT_a1_b[2]\ : OR2B
      port map(A => alu_sample(1), B => alu_coef_s(2), Y => 
        \a1_b[2]\);
    
    RESMULT_madd_126 : NOR3B
      port map(A => N_39, B => N_51, C => N_28, Y => N_56);
    
    \RESMULT_a_i14_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(14), Y => 
        \a_i14_b[8]\);
    
    RESMULT_madd_493_6 : XOR2
      port map(A => madd_493_6_0, B => N_186_1, Y => N_205);
    
    \RESMULT_a14_b[5]\ : OR2B
      port map(A => alu_sample(14), B => alu_coef_s(5), Y => 
        \a14_b[5]\);
    
    RESMULT_madd_161 : AO13
      port map(A => madd_119_m6, B => N_65_i, C => N_67, Y => 
        N_70);
    
    RESMULT_madd_606_ADD_22x22_fast_I194_Y_0_0 : XOR3
      port map(A => N_69, B => madd_124_m6, C => N_56, Y => 
        ADD_22x22_fast_I194_Y_0_0);
    
    RESMULT_madd_606_ADD_22x22_fast_I153_un1_Y : OA1A
      port map(A => I133_un1_Y_i, B => N413, C => 
        ADD_22x22_fast_I153_un1_Y_0, Y => I153_un1_Y);
    
    \RESMULT_a4_b[0]\ : OR2B
      port map(A => alu_sample(4), B => alu_coef_s(0), Y => 
        \a4_b[0]\);
    
    \RESMULT_a12_b[4]\ : OR2B
      port map(A => alu_sample(12), B => alu_coef_s(4), Y => 
        \a12_b[4]\);
    
    RESMULT_madd_205 : MAJ3
      port map(A => \a11_b[0]\, B => \a9_b[2]\, C => \a10_b[1]\, 
        Y => N_90_i);
    
    RESMULT_madd_13 : AO13
      port map(A => N_2, B => \a0_b[3]\, C => N_3, Y => N_6);
    
    RESMULT_madd_606_ADD_22x22_fast_I207_Y_0 : AX1E
      port map(A => I172_un1_Y, B => ADD_22x22_fast_I172_Y_2, C
         => ADD_22x22_fast_I207_Y_0_0, Y => \RESMULT[22]\);
    
    RESMULT_madd_606_ADD_22x22_fast_I7_G0N : NOR2B
      port map(A => N_119, B => N_104, Y => N294);
    
    RESMULT_madd_606_ADD_22x22_fast_I30_Y : AO13
      port map(A => N318, B => N_243, C => N_236, Y => N346);
    
    \RESMULT_a_i8_b[8]\ : OR2A
      port map(A => alu_coef_s(8), B => alu_sample(8), Y => 
        \a_i8_b[8]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MAC is

    port( sample_out_s : out   std_logic_vector(17 downto 0);
          alu_sample   : in    std_logic_vector(17 downto 0);
          alu_coef_s   : in    std_logic_vector(8 downto 0);
          alu_ctrl     : in    std_logic_vector(2 downto 0);
          HCLK_c       : in    std_logic;
          HRESETn_c    : in    std_logic
        );

end MAC;

architecture DEF_ARCH of MAC is 

  component MAC_REG_18
    port( alu_sample : in    std_logic_vector(17 downto 0) := (others => 'U');
          OP1_2C_D   : out   std_logic_vector(17 downto 0);
          HRESETn_c  : in    std_logic := 'U';
          HCLK_c     : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MAC_REG_9
    port( alu_coef_s : in    std_logic_vector(8 downto 0) := (others => 'U');
          OP2_2C_D   : out   std_logic_vector(8 downto 0);
          HRESETn_c  : in    std_logic := 'U';
          HCLK_c     : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component MAC_REG_1_4
    port( MACMUX2sel_D   : in    std_logic := 'U';
          HRESETn_c      : in    std_logic := 'U';
          HCLK_c         : in    std_logic := 'U';
          MACMUX2sel_D_D : out   std_logic
        );
  end component;

  component MAC_CONTROLER
    port( alu_ctrl   : in    std_logic_vector(1 downto 0) := (others => 'U');
          MACMUX2sel : out   std_logic;
          N_4        : out   std_logic;
          mult       : out   std_logic;
          mult_0     : out   std_logic
        );
  end component;

  component MAC_MUX
    port( OP1_2C_D      : in    std_logic_vector(17 downto 0) := (others => 'U');
          MULTout       : in    std_logic_vector(24 downto 0) := (others => 'U');
          ADDERinB      : out   std_logic_vector(24 downto 0);
          ADDERinA_i    : out   std_logic_vector(18 to 18);
          OP2_2C_D      : in    std_logic_vector(8 downto 0) := (others => 'U');
          ADDERout      : in    std_logic_vector(24 downto 0) := (others => 'U');
          ADDERinA_17   : out   std_logic;
          ADDERinA_24   : out   std_logic;
          ADDERinA_23   : out   std_logic;
          ADDERinA_22   : out   std_logic;
          ADDERinA_21   : out   std_logic;
          ADDERinA_20   : out   std_logic;
          ADDERinA_19   : out   std_logic;
          ADDERinA_16   : out   std_logic;
          ADDERinA_15   : out   std_logic;
          ADDERinA_14   : out   std_logic;
          ADDERinA_13   : out   std_logic;
          ADDERinA_12   : out   std_logic;
          ADDERinA_11   : out   std_logic;
          ADDERinA_10   : out   std_logic;
          ADDERinA_9    : out   std_logic;
          ADDERinA_8    : out   std_logic;
          ADDERinA_7    : out   std_logic;
          ADDERinA_6    : out   std_logic;
          ADDERinA_5    : out   std_logic;
          ADDERinA_4    : out   std_logic;
          ADDERinA_3    : out   std_logic;
          ADDERinA_2    : out   std_logic;
          ADDERinA_1    : out   std_logic;
          ADDERinA_0    : out   std_logic;
          MACMUXsel_D   : in    std_logic := 'U';
          MACMUXsel_D_1 : in    std_logic := 'U';
          MACMUXsel_D_0 : in    std_logic := 'U'
        );
  end component;

  component MAC_REG_27
    port( MULTout   : in    std_logic_vector(24 downto 7) := (others => 'U');
          MULTout_D : out   std_logic_vector(24 downto 7);
          HRESETn_c : in    std_logic := 'U';
          HCLK_c    : in    std_logic := 'U'
        );
  end component;

  component MAC_REG_1_1
    port( alu_ctrl  : in    std_logic_vector(0 to 0) := (others => 'U');
          add_D     : out   std_logic;
          HRESETn_c : in    std_logic := 'U';
          HCLK_c    : in    std_logic := 'U';
          add_D_0   : out   std_logic
        );
  end component;

  component MAC_REG_1_3
    port( MACMUX2sel   : in    std_logic := 'U';
          HRESETn_c    : in    std_logic := 'U';
          HCLK_c       : in    std_logic := 'U';
          MACMUX2sel_D : out   std_logic
        );
  end component;

  component MAC_REG_1
    port( alu_ctrl    : in    std_logic_vector(2 to 2) := (others => 'U');
          clr_MAC_D   : out   std_logic;
          HRESETn_c   : in    std_logic := 'U';
          HCLK_c      : in    std_logic := 'U';
          clr_MAC_D_0 : out   std_logic
        );
  end component;

  component Adder
    port( ADDERout     : out   std_logic_vector(24 downto 0);
          ADDERinA_i   : in    std_logic_vector(18 to 18) := (others => 'U');
          ADDERinB     : in    std_logic_vector(24 downto 0) := (others => 'U');
          ADDERinA_0   : in    std_logic := 'U';
          ADDERinA_1   : in    std_logic := 'U';
          ADDERinA_3   : in    std_logic := 'U';
          ADDERinA_5   : in    std_logic := 'U';
          ADDERinA_7   : in    std_logic := 'U';
          ADDERinA_8   : in    std_logic := 'U';
          ADDERinA_15  : in    std_logic := 'U';
          ADDERinA_16  : in    std_logic := 'U';
          ADDERinA_2   : in    std_logic := 'U';
          ADDERinA_14  : in    std_logic := 'U';
          ADDERinA_6   : in    std_logic := 'U';
          ADDERinA_10  : in    std_logic := 'U';
          ADDERinA_4   : in    std_logic := 'U';
          ADDERinA_12  : in    std_logic := 'U';
          ADDERinA_20  : in    std_logic := 'U';
          ADDERinA_11  : in    std_logic := 'U';
          ADDERinA_19  : in    std_logic := 'U';
          ADDERinA_9   : in    std_logic := 'U';
          ADDERinA_13  : in    std_logic := 'U';
          ADDERinA_21  : in    std_logic := 'U';
          ADDERinA_22  : in    std_logic := 'U';
          ADDERinA_24  : in    std_logic := 'U';
          ADDERinA_23  : in    std_logic := 'U';
          ADDERinA_17  : in    std_logic := 'U';
          HRESETn_c    : in    std_logic := 'U';
          HCLK_c       : in    std_logic := 'U';
          clr_MAC_D    : in    std_logic := 'U';
          add_D        : in    std_logic := 'U';
          clr_MAC_D_0  : in    std_logic := 'U';
          MACMUX2sel_D : in    std_logic := 'U';
          add_D_0      : in    std_logic := 'U'
        );
  end component;

  component MAC_MUX2
    port( MULTout_D      : in    std_logic_vector(24 downto 7) := (others => 'U');
          ADDERout       : in    std_logic_vector(24 downto 7) := (others => 'U');
          sample_out_s   : out   std_logic_vector(17 downto 0);
          MACMUX2sel_D_D : in    std_logic := 'U'
        );
  end component;

  component MAC_REG_1_2
    port( MACMUXsel_D   : out   std_logic;
          MACMUXsel_D_0 : out   std_logic;
          N_4           : in    std_logic := 'U';
          HRESETn_c     : in    std_logic := 'U';
          HCLK_c        : in    std_logic := 'U';
          MACMUXsel_D_1 : out   std_logic
        );
  end component;

  component Multiplier
    port( MULTout    : out   std_logic_vector(24 downto 0);
          alu_coef_s : in    std_logic_vector(8 downto 0) := (others => 'U');
          alu_sample : in    std_logic_vector(17 downto 0) := (others => 'U');
          mult       : in    std_logic := 'U';
          mult_0     : in    std_logic := 'U';
          HRESETn_c  : in    std_logic := 'U';
          HCLK_c     : in    std_logic := 'U'
        );
  end component;

    signal MACMUX2sel, N_4, mult, mult_0, \MULTout[0]\, 
        \MULTout[1]\, \MULTout[2]\, \MULTout[3]\, \MULTout[4]\, 
        \MULTout[5]\, \MULTout[6]\, \MULTout[7]\, \MULTout[8]\, 
        \MULTout[9]\, \MULTout[10]\, \MULTout[11]\, \MULTout[12]\, 
        \MULTout[13]\, \MULTout[14]\, \MULTout[15]\, 
        \MULTout[16]\, \MULTout[17]\, \MULTout[18]\, 
        \MULTout[19]\, \MULTout[20]\, \MULTout[21]\, 
        \MULTout[22]\, \MULTout[23]\, \MULTout[24]\, 
        \ADDERout[0]\, \ADDERout[1]\, \ADDERout[2]\, 
        \ADDERout[3]\, \ADDERout[4]\, \ADDERout[5]\, 
        \ADDERout[6]\, \ADDERout[7]\, \ADDERout[8]\, 
        \ADDERout[9]\, \ADDERout[10]\, \ADDERout[11]\, 
        \ADDERout[12]\, \ADDERout[13]\, \ADDERout[14]\, 
        \ADDERout[15]\, \ADDERout[16]\, \ADDERout[17]\, 
        \ADDERout[18]\, \ADDERout[19]\, \ADDERout[20]\, 
        \ADDERout[21]\, \ADDERout[22]\, \ADDERout[23]\, 
        \ADDERout[24]\, \ADDERinA_i[18]\, \ADDERinB[0]\, 
        \ADDERinB[1]\, \ADDERinB[2]\, \ADDERinB[3]\, 
        \ADDERinB[4]\, \ADDERinB[5]\, \ADDERinB[6]\, 
        \ADDERinB[7]\, \ADDERinB[8]\, \ADDERinB[9]\, 
        \ADDERinB[10]\, \ADDERinB[11]\, \ADDERinB[12]\, 
        \ADDERinB[13]\, \ADDERinB[14]\, \ADDERinB[15]\, 
        \ADDERinB[16]\, \ADDERinB[17]\, \ADDERinB[18]\, 
        \ADDERinB[19]\, \ADDERinB[20]\, \ADDERinB[21]\, 
        \ADDERinB[22]\, \ADDERinB[23]\, \ADDERinB[24]\, 
        \ADDERinA[0]\, \ADDERinA[1]\, \ADDERinA[3]\, 
        \ADDERinA[5]\, \ADDERinA[7]\, \ADDERinA[8]\, 
        \ADDERinA[15]\, \ADDERinA[16]\, \ADDERinA[2]\, 
        \ADDERinA[14]\, \ADDERinA[6]\, \ADDERinA[10]\, 
        \ADDERinA[4]\, \ADDERinA[12]\, \ADDERinA[20]\, 
        \ADDERinA[11]\, \ADDERinA[19]\, \ADDERinA[9]\, 
        \ADDERinA[13]\, \ADDERinA[21]\, \ADDERinA[22]\, 
        \ADDERinA[24]\, \ADDERinA[23]\, \ADDERinA[17]\, clr_MAC_D, 
        add_D, clr_MAC_D_0, MACMUX2sel_D, add_D_0, \OP1_2C_D[0]\, 
        \OP1_2C_D[1]\, \OP1_2C_D[2]\, \OP1_2C_D[3]\, 
        \OP1_2C_D[4]\, \OP1_2C_D[5]\, \OP1_2C_D[6]\, 
        \OP1_2C_D[7]\, \OP1_2C_D[8]\, \OP1_2C_D[9]\, 
        \OP1_2C_D[10]\, \OP1_2C_D[11]\, \OP1_2C_D[12]\, 
        \OP1_2C_D[13]\, \OP1_2C_D[14]\, \OP1_2C_D[15]\, 
        \OP1_2C_D[16]\, \OP1_2C_D[17]\, \OP2_2C_D[0]\, 
        \OP2_2C_D[1]\, \OP2_2C_D[2]\, \OP2_2C_D[3]\, 
        \OP2_2C_D[4]\, \OP2_2C_D[5]\, \OP2_2C_D[6]\, 
        \OP2_2C_D[7]\, \OP2_2C_D[8]\, \MULTout_D[7]\, 
        \MULTout_D[8]\, \MULTout_D[9]\, \MULTout_D[10]\, 
        \MULTout_D[11]\, \MULTout_D[12]\, \MULTout_D[13]\, 
        \MULTout_D[14]\, \MULTout_D[15]\, \MULTout_D[16]\, 
        \MULTout_D[17]\, \MULTout_D[18]\, \MULTout_D[19]\, 
        \MULTout_D[20]\, \MULTout_D[21]\, \MULTout_D[22]\, 
        \MULTout_D[23]\, \MULTout_D[24]\, MACMUXsel_D, 
        MACMUXsel_D_0, MACMUXsel_D_1, MACMUX2sel_D_D, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

    for all : MAC_REG_18
	Use entity work.MAC_REG_18(DEF_ARCH);
    for all : MAC_REG_9
	Use entity work.MAC_REG_9(DEF_ARCH);
    for all : MAC_REG_1_4
	Use entity work.MAC_REG_1_4(DEF_ARCH);
    for all : MAC_CONTROLER
	Use entity work.MAC_CONTROLER(DEF_ARCH);
    for all : MAC_MUX
	Use entity work.MAC_MUX(DEF_ARCH);
    for all : MAC_REG_27
	Use entity work.MAC_REG_27(DEF_ARCH);
    for all : MAC_REG_1_1
	Use entity work.MAC_REG_1_1(DEF_ARCH);
    for all : MAC_REG_1_3
	Use entity work.MAC_REG_1_3(DEF_ARCH);
    for all : MAC_REG_1
	Use entity work.MAC_REG_1(DEF_ARCH);
    for all : Adder
	Use entity work.Adder(DEF_ARCH);
    for all : MAC_MUX2
	Use entity work.MAC_MUX2(DEF_ARCH);
    for all : MAC_REG_1_2
	Use entity work.MAC_REG_1_2(DEF_ARCH);
    for all : Multiplier
	Use entity work.Multiplier(DEF_ARCH);
begin 


    OP1REG : MAC_REG_18
      port map(alu_sample(17) => alu_sample(17), alu_sample(16)
         => alu_sample(16), alu_sample(15) => alu_sample(15), 
        alu_sample(14) => alu_sample(14), alu_sample(13) => 
        alu_sample(13), alu_sample(12) => alu_sample(12), 
        alu_sample(11) => alu_sample(11), alu_sample(10) => 
        alu_sample(10), alu_sample(9) => alu_sample(9), 
        alu_sample(8) => alu_sample(8), alu_sample(7) => 
        alu_sample(7), alu_sample(6) => alu_sample(6), 
        alu_sample(5) => alu_sample(5), alu_sample(4) => 
        alu_sample(4), alu_sample(3) => alu_sample(3), 
        alu_sample(2) => alu_sample(2), alu_sample(1) => 
        alu_sample(1), alu_sample(0) => alu_sample(0), 
        OP1_2C_D(17) => \OP1_2C_D[17]\, OP1_2C_D(16) => 
        \OP1_2C_D[16]\, OP1_2C_D(15) => \OP1_2C_D[15]\, 
        OP1_2C_D(14) => \OP1_2C_D[14]\, OP1_2C_D(13) => 
        \OP1_2C_D[13]\, OP1_2C_D(12) => \OP1_2C_D[12]\, 
        OP1_2C_D(11) => \OP1_2C_D[11]\, OP1_2C_D(10) => 
        \OP1_2C_D[10]\, OP1_2C_D(9) => \OP1_2C_D[9]\, OP1_2C_D(8)
         => \OP1_2C_D[8]\, OP1_2C_D(7) => \OP1_2C_D[7]\, 
        OP1_2C_D(6) => \OP1_2C_D[6]\, OP1_2C_D(5) => 
        \OP1_2C_D[5]\, OP1_2C_D(4) => \OP1_2C_D[4]\, OP1_2C_D(3)
         => \OP1_2C_D[3]\, OP1_2C_D(2) => \OP1_2C_D[2]\, 
        OP1_2C_D(1) => \OP1_2C_D[1]\, OP1_2C_D(0) => 
        \OP1_2C_D[0]\, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    OP2REG : MAC_REG_9
      port map(alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0), 
        OP2_2C_D(8) => \OP2_2C_D[8]\, OP2_2C_D(7) => 
        \OP2_2C_D[7]\, OP2_2C_D(6) => \OP2_2C_D[6]\, OP2_2C_D(5)
         => \OP2_2C_D[5]\, OP2_2C_D(4) => \OP2_2C_D[4]\, 
        OP2_2C_D(3) => \OP2_2C_D[3]\, OP2_2C_D(2) => 
        \OP2_2C_D[2]\, OP2_2C_D(1) => \OP2_2C_D[1]\, OP2_2C_D(0)
         => \OP2_2C_D[0]\, HRESETn_c => HRESETn_c, HCLK_c => 
        HCLK_c);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    MACMUX2selREG2 : MAC_REG_1_4
      port map(MACMUX2sel_D => MACMUX2sel_D, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, MACMUX2sel_D_D => 
        MACMUX2sel_D_D);
    
    MAC_CONTROLER1 : MAC_CONTROLER
      port map(alu_ctrl(1) => alu_ctrl(1), alu_ctrl(0) => 
        alu_ctrl(0), MACMUX2sel => MACMUX2sel, N_4 => N_4, mult
         => mult, mult_0 => mult_0);
    
    MACMUX_inst : MAC_MUX
      port map(OP1_2C_D(17) => \OP1_2C_D[17]\, OP1_2C_D(16) => 
        \OP1_2C_D[16]\, OP1_2C_D(15) => \OP1_2C_D[15]\, 
        OP1_2C_D(14) => \OP1_2C_D[14]\, OP1_2C_D(13) => 
        \OP1_2C_D[13]\, OP1_2C_D(12) => \OP1_2C_D[12]\, 
        OP1_2C_D(11) => \OP1_2C_D[11]\, OP1_2C_D(10) => 
        \OP1_2C_D[10]\, OP1_2C_D(9) => \OP1_2C_D[9]\, OP1_2C_D(8)
         => \OP1_2C_D[8]\, OP1_2C_D(7) => \OP1_2C_D[7]\, 
        OP1_2C_D(6) => \OP1_2C_D[6]\, OP1_2C_D(5) => 
        \OP1_2C_D[5]\, OP1_2C_D(4) => \OP1_2C_D[4]\, OP1_2C_D(3)
         => \OP1_2C_D[3]\, OP1_2C_D(2) => \OP1_2C_D[2]\, 
        OP1_2C_D(1) => \OP1_2C_D[1]\, OP1_2C_D(0) => 
        \OP1_2C_D[0]\, MULTout(24) => \MULTout[24]\, MULTout(23)
         => \MULTout[23]\, MULTout(22) => \MULTout[22]\, 
        MULTout(21) => \MULTout[21]\, MULTout(20) => 
        \MULTout[20]\, MULTout(19) => \MULTout[19]\, MULTout(18)
         => \MULTout[18]\, MULTout(17) => \MULTout[17]\, 
        MULTout(16) => \MULTout[16]\, MULTout(15) => 
        \MULTout[15]\, MULTout(14) => \MULTout[14]\, MULTout(13)
         => \MULTout[13]\, MULTout(12) => \MULTout[12]\, 
        MULTout(11) => \MULTout[11]\, MULTout(10) => 
        \MULTout[10]\, MULTout(9) => \MULTout[9]\, MULTout(8) => 
        \MULTout[8]\, MULTout(7) => \MULTout[7]\, MULTout(6) => 
        \MULTout[6]\, MULTout(5) => \MULTout[5]\, MULTout(4) => 
        \MULTout[4]\, MULTout(3) => \MULTout[3]\, MULTout(2) => 
        \MULTout[2]\, MULTout(1) => \MULTout[1]\, MULTout(0) => 
        \MULTout[0]\, ADDERinB(24) => \ADDERinB[24]\, 
        ADDERinB(23) => \ADDERinB[23]\, ADDERinB(22) => 
        \ADDERinB[22]\, ADDERinB(21) => \ADDERinB[21]\, 
        ADDERinB(20) => \ADDERinB[20]\, ADDERinB(19) => 
        \ADDERinB[19]\, ADDERinB(18) => \ADDERinB[18]\, 
        ADDERinB(17) => \ADDERinB[17]\, ADDERinB(16) => 
        \ADDERinB[16]\, ADDERinB(15) => \ADDERinB[15]\, 
        ADDERinB(14) => \ADDERinB[14]\, ADDERinB(13) => 
        \ADDERinB[13]\, ADDERinB(12) => \ADDERinB[12]\, 
        ADDERinB(11) => \ADDERinB[11]\, ADDERinB(10) => 
        \ADDERinB[10]\, ADDERinB(9) => \ADDERinB[9]\, ADDERinB(8)
         => \ADDERinB[8]\, ADDERinB(7) => \ADDERinB[7]\, 
        ADDERinB(6) => \ADDERinB[6]\, ADDERinB(5) => 
        \ADDERinB[5]\, ADDERinB(4) => \ADDERinB[4]\, ADDERinB(3)
         => \ADDERinB[3]\, ADDERinB(2) => \ADDERinB[2]\, 
        ADDERinB(1) => \ADDERinB[1]\, ADDERinB(0) => 
        \ADDERinB[0]\, ADDERinA_i(18) => \ADDERinA_i[18]\, 
        OP2_2C_D(8) => \OP2_2C_D[8]\, OP2_2C_D(7) => 
        \OP2_2C_D[7]\, OP2_2C_D(6) => \OP2_2C_D[6]\, OP2_2C_D(5)
         => \OP2_2C_D[5]\, OP2_2C_D(4) => \OP2_2C_D[4]\, 
        OP2_2C_D(3) => \OP2_2C_D[3]\, OP2_2C_D(2) => 
        \OP2_2C_D[2]\, OP2_2C_D(1) => \OP2_2C_D[1]\, OP2_2C_D(0)
         => \OP2_2C_D[0]\, ADDERout(24) => \ADDERout[24]\, 
        ADDERout(23) => \ADDERout[23]\, ADDERout(22) => 
        \ADDERout[22]\, ADDERout(21) => \ADDERout[21]\, 
        ADDERout(20) => \ADDERout[20]\, ADDERout(19) => 
        \ADDERout[19]\, ADDERout(18) => \ADDERout[18]\, 
        ADDERout(17) => \ADDERout[17]\, ADDERout(16) => 
        \ADDERout[16]\, ADDERout(15) => \ADDERout[15]\, 
        ADDERout(14) => \ADDERout[14]\, ADDERout(13) => 
        \ADDERout[13]\, ADDERout(12) => \ADDERout[12]\, 
        ADDERout(11) => \ADDERout[11]\, ADDERout(10) => 
        \ADDERout[10]\, ADDERout(9) => \ADDERout[9]\, ADDERout(8)
         => \ADDERout[8]\, ADDERout(7) => \ADDERout[7]\, 
        ADDERout(6) => \ADDERout[6]\, ADDERout(5) => 
        \ADDERout[5]\, ADDERout(4) => \ADDERout[4]\, ADDERout(3)
         => \ADDERout[3]\, ADDERout(2) => \ADDERout[2]\, 
        ADDERout(1) => \ADDERout[1]\, ADDERout(0) => 
        \ADDERout[0]\, ADDERinA_17 => \ADDERinA[17]\, ADDERinA_24
         => \ADDERinA[24]\, ADDERinA_23 => \ADDERinA[23]\, 
        ADDERinA_22 => \ADDERinA[22]\, ADDERinA_21 => 
        \ADDERinA[21]\, ADDERinA_20 => \ADDERinA[20]\, 
        ADDERinA_19 => \ADDERinA[19]\, ADDERinA_16 => 
        \ADDERinA[16]\, ADDERinA_15 => \ADDERinA[15]\, 
        ADDERinA_14 => \ADDERinA[14]\, ADDERinA_13 => 
        \ADDERinA[13]\, ADDERinA_12 => \ADDERinA[12]\, 
        ADDERinA_11 => \ADDERinA[11]\, ADDERinA_10 => 
        \ADDERinA[10]\, ADDERinA_9 => \ADDERinA[9]\, ADDERinA_8
         => \ADDERinA[8]\, ADDERinA_7 => \ADDERinA[7]\, 
        ADDERinA_6 => \ADDERinA[6]\, ADDERinA_5 => \ADDERinA[5]\, 
        ADDERinA_4 => \ADDERinA[4]\, ADDERinA_3 => \ADDERinA[3]\, 
        ADDERinA_2 => \ADDERinA[2]\, ADDERinA_1 => \ADDERinA[1]\, 
        ADDERinA_0 => \ADDERinA[0]\, MACMUXsel_D => MACMUXsel_D, 
        MACMUXsel_D_1 => MACMUXsel_D_1, MACMUXsel_D_0 => 
        MACMUXsel_D_0);
    
    MULToutREG : MAC_REG_27
      port map(MULTout(24) => \MULTout[24]\, MULTout(23) => 
        \MULTout[23]\, MULTout(22) => \MULTout[22]\, MULTout(21)
         => \MULTout[21]\, MULTout(20) => \MULTout[20]\, 
        MULTout(19) => \MULTout[19]\, MULTout(18) => 
        \MULTout[18]\, MULTout(17) => \MULTout[17]\, MULTout(16)
         => \MULTout[16]\, MULTout(15) => \MULTout[15]\, 
        MULTout(14) => \MULTout[14]\, MULTout(13) => 
        \MULTout[13]\, MULTout(12) => \MULTout[12]\, MULTout(11)
         => \MULTout[11]\, MULTout(10) => \MULTout[10]\, 
        MULTout(9) => \MULTout[9]\, MULTout(8) => \MULTout[8]\, 
        MULTout(7) => \MULTout[7]\, MULTout_D(24) => 
        \MULTout_D[24]\, MULTout_D(23) => \MULTout_D[23]\, 
        MULTout_D(22) => \MULTout_D[22]\, MULTout_D(21) => 
        \MULTout_D[21]\, MULTout_D(20) => \MULTout_D[20]\, 
        MULTout_D(19) => \MULTout_D[19]\, MULTout_D(18) => 
        \MULTout_D[18]\, MULTout_D(17) => \MULTout_D[17]\, 
        MULTout_D(16) => \MULTout_D[16]\, MULTout_D(15) => 
        \MULTout_D[15]\, MULTout_D(14) => \MULTout_D[14]\, 
        MULTout_D(13) => \MULTout_D[13]\, MULTout_D(12) => 
        \MULTout_D[12]\, MULTout_D(11) => \MULTout_D[11]\, 
        MULTout_D(10) => \MULTout_D[10]\, MULTout_D(9) => 
        \MULTout_D[9]\, MULTout_D(8) => \MULTout_D[8]\, 
        MULTout_D(7) => \MULTout_D[7]\, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c);
    
    GND_i : GND
      port map(Y => \GND\);
    
    addREG : MAC_REG_1_1
      port map(alu_ctrl(0) => alu_ctrl(0), add_D => add_D, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, add_D_0 => 
        add_D_0);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    MACMUX2selREG : MAC_REG_1_3
      port map(MACMUX2sel => MACMUX2sel, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, MACMUX2sel_D => MACMUX2sel_D);
    
    clr_MACREG1 : MAC_REG_1
      port map(alu_ctrl(2) => alu_ctrl(2), clr_MAC_D => clr_MAC_D, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, clr_MAC_D_0 => 
        clr_MAC_D_0);
    
    adder_inst : Adder
      port map(ADDERout(24) => \ADDERout[24]\, ADDERout(23) => 
        \ADDERout[23]\, ADDERout(22) => \ADDERout[22]\, 
        ADDERout(21) => \ADDERout[21]\, ADDERout(20) => 
        \ADDERout[20]\, ADDERout(19) => \ADDERout[19]\, 
        ADDERout(18) => \ADDERout[18]\, ADDERout(17) => 
        \ADDERout[17]\, ADDERout(16) => \ADDERout[16]\, 
        ADDERout(15) => \ADDERout[15]\, ADDERout(14) => 
        \ADDERout[14]\, ADDERout(13) => \ADDERout[13]\, 
        ADDERout(12) => \ADDERout[12]\, ADDERout(11) => 
        \ADDERout[11]\, ADDERout(10) => \ADDERout[10]\, 
        ADDERout(9) => \ADDERout[9]\, ADDERout(8) => 
        \ADDERout[8]\, ADDERout(7) => \ADDERout[7]\, ADDERout(6)
         => \ADDERout[6]\, ADDERout(5) => \ADDERout[5]\, 
        ADDERout(4) => \ADDERout[4]\, ADDERout(3) => 
        \ADDERout[3]\, ADDERout(2) => \ADDERout[2]\, ADDERout(1)
         => \ADDERout[1]\, ADDERout(0) => \ADDERout[0]\, 
        ADDERinA_i(18) => \ADDERinA_i[18]\, ADDERinB(24) => 
        \ADDERinB[24]\, ADDERinB(23) => \ADDERinB[23]\, 
        ADDERinB(22) => \ADDERinB[22]\, ADDERinB(21) => 
        \ADDERinB[21]\, ADDERinB(20) => \ADDERinB[20]\, 
        ADDERinB(19) => \ADDERinB[19]\, ADDERinB(18) => 
        \ADDERinB[18]\, ADDERinB(17) => \ADDERinB[17]\, 
        ADDERinB(16) => \ADDERinB[16]\, ADDERinB(15) => 
        \ADDERinB[15]\, ADDERinB(14) => \ADDERinB[14]\, 
        ADDERinB(13) => \ADDERinB[13]\, ADDERinB(12) => 
        \ADDERinB[12]\, ADDERinB(11) => \ADDERinB[11]\, 
        ADDERinB(10) => \ADDERinB[10]\, ADDERinB(9) => 
        \ADDERinB[9]\, ADDERinB(8) => \ADDERinB[8]\, ADDERinB(7)
         => \ADDERinB[7]\, ADDERinB(6) => \ADDERinB[6]\, 
        ADDERinB(5) => \ADDERinB[5]\, ADDERinB(4) => 
        \ADDERinB[4]\, ADDERinB(3) => \ADDERinB[3]\, ADDERinB(2)
         => \ADDERinB[2]\, ADDERinB(1) => \ADDERinB[1]\, 
        ADDERinB(0) => \ADDERinB[0]\, ADDERinA_0 => \ADDERinA[0]\, 
        ADDERinA_1 => \ADDERinA[1]\, ADDERinA_3 => \ADDERinA[3]\, 
        ADDERinA_5 => \ADDERinA[5]\, ADDERinA_7 => \ADDERinA[7]\, 
        ADDERinA_8 => \ADDERinA[8]\, ADDERinA_15 => 
        \ADDERinA[15]\, ADDERinA_16 => \ADDERinA[16]\, ADDERinA_2
         => \ADDERinA[2]\, ADDERinA_14 => \ADDERinA[14]\, 
        ADDERinA_6 => \ADDERinA[6]\, ADDERinA_10 => 
        \ADDERinA[10]\, ADDERinA_4 => \ADDERinA[4]\, ADDERinA_12
         => \ADDERinA[12]\, ADDERinA_20 => \ADDERinA[20]\, 
        ADDERinA_11 => \ADDERinA[11]\, ADDERinA_19 => 
        \ADDERinA[19]\, ADDERinA_9 => \ADDERinA[9]\, ADDERinA_13
         => \ADDERinA[13]\, ADDERinA_21 => \ADDERinA[21]\, 
        ADDERinA_22 => \ADDERinA[22]\, ADDERinA_24 => 
        \ADDERinA[24]\, ADDERinA_23 => \ADDERinA[23]\, 
        ADDERinA_17 => \ADDERinA[17]\, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, clr_MAC_D => clr_MAC_D, add_D => add_D, 
        clr_MAC_D_0 => clr_MAC_D_0, MACMUX2sel_D => MACMUX2sel_D, 
        add_D_0 => add_D_0);
    
    MAC_MUX2_inst : MAC_MUX2
      port map(MULTout_D(24) => \MULTout_D[24]\, MULTout_D(23)
         => \MULTout_D[23]\, MULTout_D(22) => \MULTout_D[22]\, 
        MULTout_D(21) => \MULTout_D[21]\, MULTout_D(20) => 
        \MULTout_D[20]\, MULTout_D(19) => \MULTout_D[19]\, 
        MULTout_D(18) => \MULTout_D[18]\, MULTout_D(17) => 
        \MULTout_D[17]\, MULTout_D(16) => \MULTout_D[16]\, 
        MULTout_D(15) => \MULTout_D[15]\, MULTout_D(14) => 
        \MULTout_D[14]\, MULTout_D(13) => \MULTout_D[13]\, 
        MULTout_D(12) => \MULTout_D[12]\, MULTout_D(11) => 
        \MULTout_D[11]\, MULTout_D(10) => \MULTout_D[10]\, 
        MULTout_D(9) => \MULTout_D[9]\, MULTout_D(8) => 
        \MULTout_D[8]\, MULTout_D(7) => \MULTout_D[7]\, 
        ADDERout(24) => \ADDERout[24]\, ADDERout(23) => 
        \ADDERout[23]\, ADDERout(22) => \ADDERout[22]\, 
        ADDERout(21) => \ADDERout[21]\, ADDERout(20) => 
        \ADDERout[20]\, ADDERout(19) => \ADDERout[19]\, 
        ADDERout(18) => \ADDERout[18]\, ADDERout(17) => 
        \ADDERout[17]\, ADDERout(16) => \ADDERout[16]\, 
        ADDERout(15) => \ADDERout[15]\, ADDERout(14) => 
        \ADDERout[14]\, ADDERout(13) => \ADDERout[13]\, 
        ADDERout(12) => \ADDERout[12]\, ADDERout(11) => 
        \ADDERout[11]\, ADDERout(10) => \ADDERout[10]\, 
        ADDERout(9) => \ADDERout[9]\, ADDERout(8) => 
        \ADDERout[8]\, ADDERout(7) => \ADDERout[7]\, 
        sample_out_s(17) => sample_out_s(17), sample_out_s(16)
         => sample_out_s(16), sample_out_s(15) => 
        sample_out_s(15), sample_out_s(14) => sample_out_s(14), 
        sample_out_s(13) => sample_out_s(13), sample_out_s(12)
         => sample_out_s(12), sample_out_s(11) => 
        sample_out_s(11), sample_out_s(10) => sample_out_s(10), 
        sample_out_s(9) => sample_out_s(9), sample_out_s(8) => 
        sample_out_s(8), sample_out_s(7) => sample_out_s(7), 
        sample_out_s(6) => sample_out_s(6), sample_out_s(5) => 
        sample_out_s(5), sample_out_s(4) => sample_out_s(4), 
        sample_out_s(3) => sample_out_s(3), sample_out_s(2) => 
        sample_out_s(2), sample_out_s(1) => sample_out_s(1), 
        sample_out_s(0) => sample_out_s(0), MACMUX2sel_D_D => 
        MACMUX2sel_D_D);
    
    MACMUXselREG : MAC_REG_1_2
      port map(MACMUXsel_D => MACMUXsel_D, MACMUXsel_D_0 => 
        MACMUXsel_D_0, N_4 => N_4, HRESETn_c => HRESETn_c, HCLK_c
         => HCLK_c, MACMUXsel_D_1 => MACMUXsel_D_1);
    
    Multiplieri_nst : Multiplier
      port map(MULTout(24) => \MULTout[24]\, MULTout(23) => 
        \MULTout[23]\, MULTout(22) => \MULTout[22]\, MULTout(21)
         => \MULTout[21]\, MULTout(20) => \MULTout[20]\, 
        MULTout(19) => \MULTout[19]\, MULTout(18) => 
        \MULTout[18]\, MULTout(17) => \MULTout[17]\, MULTout(16)
         => \MULTout[16]\, MULTout(15) => \MULTout[15]\, 
        MULTout(14) => \MULTout[14]\, MULTout(13) => 
        \MULTout[13]\, MULTout(12) => \MULTout[12]\, MULTout(11)
         => \MULTout[11]\, MULTout(10) => \MULTout[10]\, 
        MULTout(9) => \MULTout[9]\, MULTout(8) => \MULTout[8]\, 
        MULTout(7) => \MULTout[7]\, MULTout(6) => \MULTout[6]\, 
        MULTout(5) => \MULTout[5]\, MULTout(4) => \MULTout[4]\, 
        MULTout(3) => \MULTout[3]\, MULTout(2) => \MULTout[2]\, 
        MULTout(1) => \MULTout[1]\, MULTout(0) => \MULTout[0]\, 
        alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0), 
        alu_sample(17) => alu_sample(17), alu_sample(16) => 
        alu_sample(16), alu_sample(15) => alu_sample(15), 
        alu_sample(14) => alu_sample(14), alu_sample(13) => 
        alu_sample(13), alu_sample(12) => alu_sample(12), 
        alu_sample(11) => alu_sample(11), alu_sample(10) => 
        alu_sample(10), alu_sample(9) => alu_sample(9), 
        alu_sample(8) => alu_sample(8), alu_sample(7) => 
        alu_sample(7), alu_sample(6) => alu_sample(6), 
        alu_sample(5) => alu_sample(5), alu_sample(4) => 
        alu_sample(4), alu_sample(3) => alu_sample(3), 
        alu_sample(2) => alu_sample(2), alu_sample(1) => 
        alu_sample(1), alu_sample(0) => alu_sample(0), mult => 
        mult, mult_0 => mult_0, HRESETn_c => HRESETn_c, HCLK_c
         => HCLK_c);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ALU is

    port( alu_ctrl     : in    std_logic_vector(2 downto 0);
          alu_coef_s   : in    std_logic_vector(8 downto 0);
          alu_sample   : in    std_logic_vector(17 downto 0);
          sample_out_s : out   std_logic_vector(17 downto 0);
          HRESETn_c    : in    std_logic;
          HCLK_c       : in    std_logic
        );

end ALU;

architecture DEF_ARCH of ALU is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MAC
    port( sample_out_s : out   std_logic_vector(17 downto 0);
          alu_sample   : in    std_logic_vector(17 downto 0) := (others => 'U');
          alu_coef_s   : in    std_logic_vector(8 downto 0) := (others => 'U');
          alu_ctrl     : in    std_logic_vector(2 downto 0) := (others => 'U');
          HCLK_c       : in    std_logic := 'U';
          HRESETn_c    : in    std_logic := 'U'
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : MAC
	Use entity work.MAC(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \arith.MACinst\ : MAC
      port map(sample_out_s(17) => sample_out_s(17), 
        sample_out_s(16) => sample_out_s(16), sample_out_s(15)
         => sample_out_s(15), sample_out_s(14) => 
        sample_out_s(14), sample_out_s(13) => sample_out_s(13), 
        sample_out_s(12) => sample_out_s(12), sample_out_s(11)
         => sample_out_s(11), sample_out_s(10) => 
        sample_out_s(10), sample_out_s(9) => sample_out_s(9), 
        sample_out_s(8) => sample_out_s(8), sample_out_s(7) => 
        sample_out_s(7), sample_out_s(6) => sample_out_s(6), 
        sample_out_s(5) => sample_out_s(5), sample_out_s(4) => 
        sample_out_s(4), sample_out_s(3) => sample_out_s(3), 
        sample_out_s(2) => sample_out_s(2), sample_out_s(1) => 
        sample_out_s(1), sample_out_s(0) => sample_out_s(0), 
        alu_sample(17) => alu_sample(17), alu_sample(16) => 
        alu_sample(16), alu_sample(15) => alu_sample(15), 
        alu_sample(14) => alu_sample(14), alu_sample(13) => 
        alu_sample(13), alu_sample(12) => alu_sample(12), 
        alu_sample(11) => alu_sample(11), alu_sample(10) => 
        alu_sample(10), alu_sample(9) => alu_sample(9), 
        alu_sample(8) => alu_sample(8), alu_sample(7) => 
        alu_sample(7), alu_sample(6) => alu_sample(6), 
        alu_sample(5) => alu_sample(5), alu_sample(4) => 
        alu_sample(4), alu_sample(3) => alu_sample(3), 
        alu_sample(2) => alu_sample(2), alu_sample(1) => 
        alu_sample(1), alu_sample(0) => alu_sample(0), 
        alu_coef_s(8) => alu_coef_s(8), alu_coef_s(7) => 
        alu_coef_s(7), alu_coef_s(6) => alu_coef_s(6), 
        alu_coef_s(5) => alu_coef_s(5), alu_coef_s(4) => 
        alu_coef_s(4), alu_coef_s(3) => alu_coef_s(3), 
        alu_coef_s(2) => alu_coef_s(2), alu_coef_s(1) => 
        alu_coef_s(1), alu_coef_s(0) => alu_coef_s(0), 
        alu_ctrl(2) => alu_ctrl(2), alu_ctrl(1) => alu_ctrl(1), 
        alu_ctrl(0) => alu_ctrl(0), HCLK_c => HCLK_c, HRESETn_c
         => HRESETn_c);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity generic_syncram_2p_8_18_0 is

    port( ram_input                     : in    std_logic_vector(17 downto 0);
          counter                       : in    std_logic_vector(7 downto 0);
          DIN_REG1_15                   : out   std_logic;
          ram_output_16                 : out   std_logic;
          ram_output_0                  : out   std_logic;
          ram_output_17                 : out   std_logic;
          ram_output_15                 : out   std_logic;
          ram_output_14                 : out   std_logic;
          ram_output_13                 : out   std_logic;
          ram_output_12                 : out   std_logic;
          ram_output_11                 : out   std_logic;
          ram_output_10                 : out   std_logic;
          ram_output_9                  : out   std_logic;
          ram_output_8                  : out   std_logic;
          ram_output_7                  : out   std_logic;
          ram_output_6                  : out   std_logic;
          ram_output_5                  : out   std_logic;
          ram_output_4                  : out   std_logic;
          ram_output_3                  : out   std_logic;
          ram_output_1                  : out   std_logic;
          reg_sample_in                 : in    std_logic_vector(6 downto 5);
          reg_sample_in_RNIFA3C         : in    std_logic_vector(15 to 15);
          alu_sample_1                  : out   std_logic;
          alu_sample_0                  : out   std_logic;
          alu_sample_10                 : out   std_logic;
          ram_write_i                   : in    std_logic;
          generic_syncram_2p_8_18_0_VCC : in    std_logic;
          generic_syncram_2p_8_18_0_GND : in    std_logic;
          ADD_8x8_medium_area_I30_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I29_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I28_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I27_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I26_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I25_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I24_Y_0   : in    std_logic;
          ADD_8x8_medium_area_I0_S_0    : in    std_logic;
          ram_write                     : in    std_logic;
          HCLK_c                        : in    std_logic;
          alu_sel_input                 : in    std_logic;
          I_1_RNI3I3E3                  : out   std_logic
        );

end generic_syncram_2p_8_18_0;

architecture DEF_ARCH of generic_syncram_2p_8_18_0 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM512X18
    generic (MEMORYFILE:string := "");

    port( RADDR8 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          WADDR8 : in    std_logic := 'U';
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          WD17   : in    std_logic := 'U';
          WD16   : in    std_logic := 'U';
          WD15   : in    std_logic := 'U';
          WD14   : in    std_logic := 'U';
          WD13   : in    std_logic := 'U';
          WD12   : in    std_logic := 'U';
          WD11   : in    std_logic := 'U';
          WD10   : in    std_logic := 'U';
          WD9    : in    std_logic := 'U';
          WD8    : in    std_logic := 'U';
          WD7    : in    std_logic := 'U';
          WD6    : in    std_logic := 'U';
          WD5    : in    std_logic := 'U';
          WD4    : in    std_logic := 'U';
          WD3    : in    std_logic := 'U';
          WD2    : in    std_logic := 'U';
          WD1    : in    std_logic := 'U';
          WD0    : in    std_logic := 'U';
          RW0    : in    std_logic := 'U';
          RW1    : in    std_logic := 'U';
          WW0    : in    std_logic := 'U';
          WW1    : in    std_logic := 'U';
          PIPE   : in    std_logic := 'U';
          REN    : in    std_logic := 'U';
          WEN    : in    std_logic := 'U';
          RCLK   : in    std_logic := 'U';
          WCLK   : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          RD17   : out   std_logic;
          RD16   : out   std_logic;
          RD15   : out   std_logic;
          RD14   : out   std_logic;
          RD13   : out   std_logic;
          RD12   : out   std_logic;
          RD11   : out   std_logic;
          RD10   : out   std_logic;
          RD9    : out   std_logic;
          RD8    : out   std_logic;
          RD7    : out   std_logic;
          RD6    : out   std_logic;
          RD5    : out   std_logic;
          RD4    : out   std_logic;
          RD3    : out   std_logic;
          RD2    : out   std_logic;
          RD1    : out   std_logic;
          RD0    : out   std_logic
        );
  end component;

    signal I_5_1, I_4_0_i_0, I_4_1_i_0, I_4_3, I_5_0, 
        \RADDR_REG1[2]\, \WADDR_REG1[2]\, N_5, I_5_2, I_5_5_0, 
        I_5_5_1, \RADDR_REG1[6]\, \WADDR_REG1[6]\, I_4_7_i_0, 
        \RADDR_REG1[4]\, \WADDR_REG1[4]\, I_4_5_i_0, N_7_i_0, 
        \DIN_REG1[2]\, \DOUT_TMP[2]\, \DOUT_TMP[15]\, 
        I_3_RNI91FA3, \DOUT_TMP[5]\, \DIN_REG1_RNIVQEG[5]\, 
        \DIN_REG1[5]\, \DOUT_TMP[6]\, \DIN_REG1_RNI13FG[6]\, 
        \DIN_REG1[6]\, \WADDR_REG1[0]\, \RADDR_REG1[0]\, 
        \WADDR_REG1[1]\, \RADDR_REG1[1]\, \WADDR_REG1[3]\, 
        \RADDR_REG1[3]\, \WADDR_REG1[5]\, \RADDR_REG1[5]\, 
        \WADDR_REG1[7]\, \RADDR_REG1[7]\, \DIN_REG1[1]\, 
        \DOUT_TMP[1]\, \DIN_REG1[3]\, \DOUT_TMP[3]\, 
        \DIN_REG1[4]\, \DOUT_TMP[4]\, \DIN_REG1[7]\, 
        \DOUT_TMP[7]\, \DIN_REG1[8]\, \DOUT_TMP[8]\, 
        \DIN_REG1[9]\, \DOUT_TMP[9]\, \DIN_REG1[10]\, 
        \DOUT_TMP[10]\, \DIN_REG1[11]\, \DOUT_TMP[11]\, 
        \DIN_REG1[12]\, \DOUT_TMP[12]\, \DIN_REG1[13]\, 
        \DOUT_TMP[13]\, \DIN_REG1[14]\, \DOUT_TMP[14]\, 
        \DIN_REG1[17]\, \DOUT_TMP[17]\, \DIN_REG1[0]\, 
        \DOUT_TMP[0]\, \DIN_REG1[16]\, \DOUT_TMP[16]\, 
        \DIN_REG1[15]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    DIN_REG1_15 <= \DIN_REG1[15]\;

    rfd_tile_I_1_RNIAE4E3 : MX2
      port map(A => \DIN_REG1[9]\, B => \DOUT_TMP[9]\, S => 
        N_7_i_0, Y => ram_output_9);
    
    rfd_tile_I_1_RNI038F3 : MX2
      port map(A => \DIN_REG1[12]\, B => \DOUT_TMP[12]\, S => 
        N_7_i_0, Y => ram_output_12);
    
    \rfd_tile_DIN_REG1_RNI13FG[6]\ : MX2
      port map(A => reg_sample_in(6), B => \DIN_REG1[6]\, S => 
        alu_sel_input, Y => \DIN_REG1_RNI13FG[6]\);
    
    \rfd_tile_DIN_REG1[9]\ : DFN1
      port map(D => ram_input(9), CLK => HCLK_c, Q => 
        \DIN_REG1[9]\);
    
    rfd_tile_I_1_RNI4M3E3 : MX2
      port map(A => \DIN_REG1[3]\, B => \DOUT_TMP[3]\, S => 
        N_7_i_0, Y => ram_output_3);
    
    \rfd_tile_RADDR_REG1[5]\ : DFN1
      port map(D => counter(5), CLK => HCLK_c, Q => 
        \RADDR_REG1[5]\);
    
    \rfd_tile_WADDR_REG1[6]\ : DFN1
      port map(D => ADD_8x8_medium_area_I29_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[6]\);
    
    rfd_tile_I_3 : DFN1
      port map(D => ram_write, CLK => HCLK_c, Q => N_5);
    
    rfd_tile_I_1_RNI2E3E3 : MX2
      port map(A => \DIN_REG1[1]\, B => \DOUT_TMP[1]\, S => 
        N_7_i_0, Y => ram_output_1);
    
    rfd_tile_I_1_RNI5Q3E3 : MX2
      port map(A => \DIN_REG1[4]\, B => \DOUT_TMP[4]\, S => 
        N_7_i_0, Y => ram_output_4);
    
    \rfd_tile_DIN_REG1[10]\ : DFN1
      port map(D => ram_input(10), CLK => HCLK_c, Q => 
        \DIN_REG1[10]\);
    
    \rfd_tile_WADDR_REG1[4]\ : DFN1
      port map(D => ADD_8x8_medium_area_I27_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[4]\);
    
    \rfd_tile_RADDR_REG1_RNIL9AC[1]\ : XNOR2
      port map(A => \WADDR_REG1[1]\, B => \RADDR_REG1[1]\, Y => 
        I_4_1_i_0);
    
    rfd_tile_I_1_RNI1A3E3 : MX2
      port map(A => \DIN_REG1[0]\, B => \DOUT_TMP[0]\, S => 
        N_7_i_0, Y => ram_output_0);
    
    rfd_tile_I_3_RNI91FA3 : OR2B
      port map(A => alu_sel_input, B => N_7_i_0, Y => 
        I_3_RNI91FA3);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \rfd_tile_DIN_REG1[0]\ : DFN1
      port map(D => ram_input(0), CLK => HCLK_c, Q => 
        \DIN_REG1[0]\);
    
    \rfd_tile_DIN_REG1[5]\ : DFN1
      port map(D => ram_input(5), CLK => HCLK_c, Q => 
        \DIN_REG1[5]\);
    
    \rfd_tile_DIN_REG1[4]\ : DFN1
      port map(D => ram_input(4), CLK => HCLK_c, Q => 
        \DIN_REG1[4]\);
    
    \rfd_tile_DIN_REG1[3]\ : DFN1
      port map(D => ram_input(3), CLK => HCLK_c, Q => 
        \DIN_REG1[3]\);
    
    \rfd_tile_DIN_REG1[2]\ : DFN1
      port map(D => ram_input(2), CLK => HCLK_c, Q => 
        \DIN_REG1[2]\);
    
    \rfd_tile_DIN_REG1[12]\ : DFN1
      port map(D => ram_input(12), CLK => HCLK_c, Q => 
        \DIN_REG1[12]\);
    
    \rfd_tile_WADDR_REG1[7]\ : DFN1
      port map(D => ADD_8x8_medium_area_I30_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[7]\);
    
    rfd_tile_I_3_RNIVS763 : OR2B
      port map(A => I_5_2, B => I_5_1, Y => N_7_i_0);
    
    rfd_tile_I_3_RNI60RF : XA1A
      port map(A => \RADDR_REG1[2]\, B => \WADDR_REG1[2]\, C => 
        N_5, Y => I_5_0);
    
    rfd_tile_I_1_RNI864E3 : MX2
      port map(A => \DIN_REG1[7]\, B => \DOUT_TMP[7]\, S => 
        N_7_i_0, Y => ram_output_7);
    
    \rfd_tile_RADDR_REG1_RNIOBMO[4]\ : XA1A
      port map(A => \RADDR_REG1[4]\, B => \WADDR_REG1[4]\, C => 
        I_4_5_i_0, Y => I_5_5_0);
    
    rfd_tile_I_1_RNIV28F3 : MX2
      port map(A => \DIN_REG1[11]\, B => \DOUT_TMP[11]\, S => 
        N_7_i_0, Y => ram_output_11);
    
    \rfd_tile_DIN_REG1[15]\ : DFN1
      port map(D => ram_input(15), CLK => HCLK_c, Q => 
        \DIN_REG1[15]\);
    
    \rfd_tile_RADDR_REG1[0]\ : DFN1
      port map(D => counter(0), CLK => HCLK_c, Q => 
        \RADDR_REG1[0]\);
    
    \rfd_tile_WADDR_REG1[5]\ : DFN1
      port map(D => ADD_8x8_medium_area_I28_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[5]\);
    
    rfd_tile_I_1_RNINIEU3 : MX2
      port map(A => \DOUT_TMP[6]\, B => \DIN_REG1_RNI13FG[6]\, S
         => I_3_RNI91FA3, Y => alu_sample_1);
    
    rfd_tile_I_1_RNI3I3E3 : MX2
      port map(A => \DIN_REG1[2]\, B => \DOUT_TMP[2]\, S => 
        N_7_i_0, Y => I_1_RNI3I3E3);
    
    \rfd_tile_RADDR_REG1[2]\ : DFN1
      port map(D => counter(2), CLK => HCLK_c, Q => 
        \RADDR_REG1[2]\);
    
    \rfd_tile_DIN_REG1[1]\ : DFN1
      port map(D => ram_input(1), CLK => HCLK_c, Q => 
        \DIN_REG1[1]\);
    
    rfd_tile_I_1_RNI5Q2Q3 : MX2
      port map(A => \DOUT_TMP[15]\, B => 
        reg_sample_in_RNIFA3C(15), S => I_3_RNI91FA3, Y => 
        alu_sample_10);
    
    \rfd_tile_RADDR_REG1[3]\ : DFN1
      port map(D => counter(3), CLK => HCLK_c, Q => 
        \RADDR_REG1[3]\);
    
    rfd_tile_I_3_RNIUN812 : NOR3C
      port map(A => I_5_5_0, B => I_5_5_1, C => I_5_0, Y => I_5_2);
    
    GND_i : GND
      port map(Y => \GND\);
    
    rfd_tile_I_1_RNI338F3 : MX2
      port map(A => \DIN_REG1[15]\, B => \DOUT_TMP[15]\, S => 
        N_7_i_0, Y => ram_output_15);
    
    \rfd_tile_RADDR_REG1_RNIT9BC[5]\ : XNOR2
      port map(A => \WADDR_REG1[5]\, B => \RADDR_REG1[5]\, Y => 
        I_4_5_i_0);
    
    \rfd_tile_RADDR_REG1[1]\ : DFN1
      port map(D => counter(1), CLK => HCLK_c, Q => 
        \RADDR_REG1[1]\);
    
    \rfd_tile_DIN_REG1_RNIVQEG[5]\ : MX2
      port map(A => reg_sample_in(5), B => \DIN_REG1[5]\, S => 
        alu_sel_input, Y => \DIN_REG1_RNIVQEG[5]\);
    
    rfd_tile_I_1_RNI9A4E3 : MX2
      port map(A => \DIN_REG1[8]\, B => \DOUT_TMP[8]\, S => 
        N_7_i_0, Y => ram_output_8);
    
    \rfd_tile_DIN_REG1[14]\ : DFN1
      port map(D => ram_input(14), CLK => HCLK_c, Q => 
        \DIN_REG1[14]\);
    
    \rfd_tile_RADDR_REG1_RNI15V41[0]\ : NOR3B
      port map(A => I_4_0_i_0, B => I_4_1_i_0, C => I_4_3, Y => 
        I_5_1);
    
    \rfd_tile_RADDR_REG1_RNIJ1AC[0]\ : XNOR2
      port map(A => \WADDR_REG1[0]\, B => \RADDR_REG1[0]\, Y => 
        I_4_0_i_0);
    
    rfd_tile_I_1_RNIU28F3 : MX2
      port map(A => \DIN_REG1[10]\, B => \DOUT_TMP[10]\, S => 
        N_7_i_0, Y => ram_output_10);
    
    \rfd_tile_RADDR_REG1[6]\ : DFN1
      port map(D => counter(6), CLK => HCLK_c, Q => 
        \RADDR_REG1[6]\);
    
    rfd_tile_I_1_RNI724E3 : MX2C
      port map(A => \DIN_REG1[6]\, B => \DOUT_TMP[6]\, S => 
        N_7_i_0, Y => ram_output_6);
    
    \rfd_tile_RADDR_REG1_RNI1QBC[7]\ : XNOR2
      port map(A => \WADDR_REG1[7]\, B => \RADDR_REG1[7]\, Y => 
        I_4_7_i_0);
    
    \rfd_tile_RADDR_REG1_RNIPPAC[3]\ : XOR2
      port map(A => \WADDR_REG1[3]\, B => \RADDR_REG1[3]\, Y => 
        I_4_3);
    
    \rfd_tile_DIN_REG1[8]\ : DFN1
      port map(D => ram_input(8), CLK => HCLK_c, Q => 
        \DIN_REG1[8]\);
    
    \rfd_tile_WADDR_REG1[0]\ : DFN1
      port map(D => ADD_8x8_medium_area_I0_S_0, CLK => HCLK_c, Q
         => \WADDR_REG1[0]\);
    
    \rfd_tile_RADDR_REG1[4]\ : DFN1
      port map(D => counter(4), CLK => HCLK_c, Q => 
        \RADDR_REG1[4]\);
    
    rfd_tile_I_1_RNI138F3 : MX2
      port map(A => \DIN_REG1[13]\, B => \DOUT_TMP[13]\, S => 
        N_7_i_0, Y => ram_output_13);
    
    \rfd_tile_DIN_REG1[6]\ : DFN1
      port map(D => ram_input(6), CLK => HCLK_c, Q => 
        \DIN_REG1[6]\);
    
    \rfd_tile_WADDR_REG1[2]\ : DFN1
      port map(D => ADD_8x8_medium_area_I25_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[2]\);
    
    \rfd_tile_DIN_REG1[11]\ : DFN1
      port map(D => ram_input(11), CLK => HCLK_c, Q => 
        \DIN_REG1[11]\);
    
    rfd_tile_I_1_RNILAEU3 : MX2
      port map(A => \DOUT_TMP[5]\, B => \DIN_REG1_RNIVQEG[5]\, S
         => I_3_RNI91FA3, Y => alu_sample_0);
    
    \rfd_tile_WADDR_REG1[3]\ : DFN1
      port map(D => ADD_8x8_medium_area_I26_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[3]\);
    
    rfd_tile_I_1_RNI438F3 : MX2
      port map(A => \DIN_REG1[16]\, B => \DOUT_TMP[16]\, S => 
        N_7_i_0, Y => ram_output_16);
    
    rfd_tile_I_1_RNI238F3 : MX2
      port map(A => \DIN_REG1[14]\, B => \DOUT_TMP[14]\, S => 
        N_7_i_0, Y => ram_output_14);
    
    \rfd_tile_DIN_REG1[13]\ : DFN1
      port map(D => ram_input(13), CLK => HCLK_c, Q => 
        \DIN_REG1[13]\);
    
    \rfd_tile_RADDR_REG1_RNI0CNO[6]\ : XA1A
      port map(A => \RADDR_REG1[6]\, B => \WADDR_REG1[6]\, C => 
        I_4_7_i_0, Y => I_5_5_1);
    
    rfd_tile_I_1_RNI538F3 : MX2
      port map(A => \DIN_REG1[17]\, B => \DOUT_TMP[17]\, S => 
        N_7_i_0, Y => ram_output_17);
    
    rfd_tile_I_1 : RAM512X18
      port map(RADDR8 => generic_syncram_2p_8_18_0_GND, RADDR7
         => counter(7), RADDR6 => counter(6), RADDR5 => 
        counter(5), RADDR4 => counter(4), RADDR3 => counter(3), 
        RADDR2 => counter(2), RADDR1 => counter(1), RADDR0 => 
        counter(0), WADDR8 => generic_syncram_2p_8_18_0_GND, 
        WADDR7 => ADD_8x8_medium_area_I30_Y_0, WADDR6 => 
        ADD_8x8_medium_area_I29_Y_0, WADDR5 => 
        ADD_8x8_medium_area_I28_Y_0, WADDR4 => 
        ADD_8x8_medium_area_I27_Y_0, WADDR3 => 
        ADD_8x8_medium_area_I26_Y_0, WADDR2 => 
        ADD_8x8_medium_area_I25_Y_0, WADDR1 => 
        ADD_8x8_medium_area_I24_Y_0, WADDR0 => 
        ADD_8x8_medium_area_I0_S_0, WD17 => ram_input(17), WD16
         => ram_input(16), WD15 => ram_input(15), WD14 => 
        ram_input(14), WD13 => ram_input(13), WD12 => 
        ram_input(12), WD11 => ram_input(11), WD10 => 
        ram_input(10), WD9 => ram_input(9), WD8 => ram_input(8), 
        WD7 => ram_input(7), WD6 => ram_input(6), WD5 => 
        ram_input(5), WD4 => ram_input(4), WD3 => ram_input(3), 
        WD2 => ram_input(2), WD1 => ram_input(1), WD0 => 
        ram_input(0), RW0 => generic_syncram_2p_8_18_0_GND, RW1
         => generic_syncram_2p_8_18_0_VCC, WW0 => 
        generic_syncram_2p_8_18_0_GND, WW1 => 
        generic_syncram_2p_8_18_0_VCC, PIPE => 
        generic_syncram_2p_8_18_0_GND, REN => 
        generic_syncram_2p_8_18_0_GND, WEN => ram_write_i, RCLK
         => HCLK_c, WCLK => HCLK_c, RESET => 
        generic_syncram_2p_8_18_0_VCC, RD17 => \DOUT_TMP[17]\, 
        RD16 => \DOUT_TMP[16]\, RD15 => \DOUT_TMP[15]\, RD14 => 
        \DOUT_TMP[14]\, RD13 => \DOUT_TMP[13]\, RD12 => 
        \DOUT_TMP[12]\, RD11 => \DOUT_TMP[11]\, RD10 => 
        \DOUT_TMP[10]\, RD9 => \DOUT_TMP[9]\, RD8 => 
        \DOUT_TMP[8]\, RD7 => \DOUT_TMP[7]\, RD6 => \DOUT_TMP[6]\, 
        RD5 => \DOUT_TMP[5]\, RD4 => \DOUT_TMP[4]\, RD3 => 
        \DOUT_TMP[3]\, RD2 => \DOUT_TMP[2]\, RD1 => \DOUT_TMP[1]\, 
        RD0 => \DOUT_TMP[0]\);
    
    \rfd_tile_RADDR_REG1[7]\ : DFN1
      port map(D => counter(7), CLK => HCLK_c, Q => 
        \RADDR_REG1[7]\);
    
    \rfd_tile_DIN_REG1[16]\ : DFN1
      port map(D => ram_input(16), CLK => HCLK_c, Q => 
        \DIN_REG1[16]\);
    
    \rfd_tile_WADDR_REG1[1]\ : DFN1
      port map(D => ADD_8x8_medium_area_I24_Y_0, CLK => HCLK_c, Q
         => \WADDR_REG1[1]\);
    
    rfd_tile_I_1_RNI6U3E3 : MX2C
      port map(A => \DIN_REG1[5]\, B => \DOUT_TMP[5]\, S => 
        N_7_i_0, Y => ram_output_5);
    
    \rfd_tile_DIN_REG1[17]\ : DFN1
      port map(D => ram_input(17), CLK => HCLK_c, Q => 
        \DIN_REG1[17]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \rfd_tile_DIN_REG1[7]\ : DFN1
      port map(D => ram_input(7), CLK => HCLK_c, Q => 
        \DIN_REG1[7]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity syncram_2pZ0 is

    port( alu_sample_10               : out   std_logic;
          alu_sample_0                : out   std_logic;
          alu_sample_1                : out   std_logic;
          reg_sample_in_RNIFA3C       : in    std_logic_vector(15 to 15);
          reg_sample_in               : in    std_logic_vector(6 downto 5);
          ram_output_1                : out   std_logic;
          ram_output_3                : out   std_logic;
          ram_output_4                : out   std_logic;
          ram_output_5                : out   std_logic;
          ram_output_6                : out   std_logic;
          ram_output_7                : out   std_logic;
          ram_output_8                : out   std_logic;
          ram_output_9                : out   std_logic;
          ram_output_10               : out   std_logic;
          ram_output_11               : out   std_logic;
          ram_output_12               : out   std_logic;
          ram_output_13               : out   std_logic;
          ram_output_14               : out   std_logic;
          ram_output_15               : out   std_logic;
          ram_output_17               : out   std_logic;
          ram_output_0                : out   std_logic;
          ram_output_16               : out   std_logic;
          DIN_REG1                    : out   std_logic_vector(15 to 15);
          counter                     : in    std_logic_vector(7 downto 0);
          ram_input                   : in    std_logic_vector(17 downto 0);
          I_1_RNI3I3E3                : out   std_logic;
          alu_sel_input               : in    std_logic;
          HCLK_c                      : in    std_logic;
          ram_write                   : in    std_logic;
          ADD_8x8_medium_area_I0_S_0  : in    std_logic;
          ADD_8x8_medium_area_I24_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I25_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I26_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I27_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I28_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I29_Y_0 : in    std_logic;
          ADD_8x8_medium_area_I30_Y_0 : in    std_logic;
          syncram_2pZ0_GND            : in    std_logic;
          syncram_2pZ0_VCC            : in    std_logic;
          ram_write_i                 : in    std_logic
        );

end syncram_2pZ0;

architecture DEF_ARCH of syncram_2pZ0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component generic_syncram_2p_8_18_0
    port( ram_input                     : in    std_logic_vector(17 downto 0) := (others => 'U');
          counter                       : in    std_logic_vector(7 downto 0) := (others => 'U');
          DIN_REG1_15                   : out   std_logic;
          ram_output_16                 : out   std_logic;
          ram_output_0                  : out   std_logic;
          ram_output_17                 : out   std_logic;
          ram_output_15                 : out   std_logic;
          ram_output_14                 : out   std_logic;
          ram_output_13                 : out   std_logic;
          ram_output_12                 : out   std_logic;
          ram_output_11                 : out   std_logic;
          ram_output_10                 : out   std_logic;
          ram_output_9                  : out   std_logic;
          ram_output_8                  : out   std_logic;
          ram_output_7                  : out   std_logic;
          ram_output_6                  : out   std_logic;
          ram_output_5                  : out   std_logic;
          ram_output_4                  : out   std_logic;
          ram_output_3                  : out   std_logic;
          ram_output_1                  : out   std_logic;
          reg_sample_in                 : in    std_logic_vector(6 downto 5) := (others => 'U');
          reg_sample_in_RNIFA3C         : in    std_logic_vector(15 to 15) := (others => 'U');
          alu_sample_1                  : out   std_logic;
          alu_sample_0                  : out   std_logic;
          alu_sample_10                 : out   std_logic;
          ram_write_i                   : in    std_logic := 'U';
          generic_syncram_2p_8_18_0_VCC : in    std_logic := 'U';
          generic_syncram_2p_8_18_0_GND : in    std_logic := 'U';
          ADD_8x8_medium_area_I30_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I29_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I28_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I27_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I26_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I25_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I24_Y_0   : in    std_logic := 'U';
          ADD_8x8_medium_area_I0_S_0    : in    std_logic := 'U';
          ram_write                     : in    std_logic := 'U';
          HCLK_c                        : in    std_logic := 'U';
          alu_sel_input                 : in    std_logic := 'U';
          I_1_RNI3I3E3                  : out   std_logic
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : generic_syncram_2p_8_18_0
	Use entity work.generic_syncram_2p_8_18_0(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \inf.x0\ : generic_syncram_2p_8_18_0
      port map(ram_input(17) => ram_input(17), ram_input(16) => 
        ram_input(16), ram_input(15) => ram_input(15), 
        ram_input(14) => ram_input(14), ram_input(13) => 
        ram_input(13), ram_input(12) => ram_input(12), 
        ram_input(11) => ram_input(11), ram_input(10) => 
        ram_input(10), ram_input(9) => ram_input(9), ram_input(8)
         => ram_input(8), ram_input(7) => ram_input(7), 
        ram_input(6) => ram_input(6), ram_input(5) => 
        ram_input(5), ram_input(4) => ram_input(4), ram_input(3)
         => ram_input(3), ram_input(2) => ram_input(2), 
        ram_input(1) => ram_input(1), ram_input(0) => 
        ram_input(0), counter(7) => counter(7), counter(6) => 
        counter(6), counter(5) => counter(5), counter(4) => 
        counter(4), counter(3) => counter(3), counter(2) => 
        counter(2), counter(1) => counter(1), counter(0) => 
        counter(0), DIN_REG1_15 => DIN_REG1(15), ram_output_16
         => ram_output_16, ram_output_0 => ram_output_0, 
        ram_output_17 => ram_output_17, ram_output_15 => 
        ram_output_15, ram_output_14 => ram_output_14, 
        ram_output_13 => ram_output_13, ram_output_12 => 
        ram_output_12, ram_output_11 => ram_output_11, 
        ram_output_10 => ram_output_10, ram_output_9 => 
        ram_output_9, ram_output_8 => ram_output_8, ram_output_7
         => ram_output_7, ram_output_6 => ram_output_6, 
        ram_output_5 => ram_output_5, ram_output_4 => 
        ram_output_4, ram_output_3 => ram_output_3, ram_output_1
         => ram_output_1, reg_sample_in(6) => reg_sample_in(6), 
        reg_sample_in(5) => reg_sample_in(5), 
        reg_sample_in_RNIFA3C(15) => reg_sample_in_RNIFA3C(15), 
        alu_sample_1 => alu_sample_1, alu_sample_0 => 
        alu_sample_0, alu_sample_10 => alu_sample_10, ram_write_i
         => ram_write_i, generic_syncram_2p_8_18_0_VCC => 
        syncram_2pZ0_VCC, generic_syncram_2p_8_18_0_GND => 
        syncram_2pZ0_GND, ADD_8x8_medium_area_I30_Y_0 => 
        ADD_8x8_medium_area_I30_Y_0, ADD_8x8_medium_area_I29_Y_0
         => ADD_8x8_medium_area_I29_Y_0, 
        ADD_8x8_medium_area_I28_Y_0 => 
        ADD_8x8_medium_area_I28_Y_0, ADD_8x8_medium_area_I27_Y_0
         => ADD_8x8_medium_area_I27_Y_0, 
        ADD_8x8_medium_area_I26_Y_0 => 
        ADD_8x8_medium_area_I26_Y_0, ADD_8x8_medium_area_I25_Y_0
         => ADD_8x8_medium_area_I25_Y_0, 
        ADD_8x8_medium_area_I24_Y_0 => 
        ADD_8x8_medium_area_I24_Y_0, ADD_8x8_medium_area_I0_S_0
         => ADD_8x8_medium_area_I0_S_0, ram_write => ram_write, 
        HCLK_c => HCLK_c, alu_sel_input => alu_sel_input, 
        I_1_RNI3I3E3 => I_1_RNI3I3E3);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity RAM_CTRLR_v2 is

    port( ram_input             : in    std_logic_vector(17 downto 0);
          DIN_REG1              : out   std_logic_vector(15 to 15);
          ram_output_16         : out   std_logic;
          ram_output_0          : out   std_logic;
          ram_output_17         : out   std_logic;
          ram_output_15         : out   std_logic;
          ram_output_14         : out   std_logic;
          ram_output_13         : out   std_logic;
          ram_output_12         : out   std_logic;
          ram_output_11         : out   std_logic;
          ram_output_10         : out   std_logic;
          ram_output_9          : out   std_logic;
          ram_output_8          : out   std_logic;
          ram_output_7          : out   std_logic;
          ram_output_6          : out   std_logic;
          ram_output_5          : out   std_logic;
          ram_output_4          : out   std_logic;
          ram_output_3          : out   std_logic;
          ram_output_1          : out   std_logic;
          reg_sample_in         : in    std_logic_vector(6 downto 5);
          reg_sample_in_RNIFA3C : in    std_logic_vector(15 to 15);
          alu_sample_1          : out   std_logic;
          alu_sample_0          : out   std_logic;
          alu_sample_10         : out   std_logic;
          waddr_previous        : in    std_logic_vector(1 downto 0);
          ram_write_i           : in    std_logic;
          RAM_CTRLR_v2_VCC      : in    std_logic;
          RAM_CTRLR_v2_GND      : in    std_logic;
          ram_write             : in    std_logic;
          alu_sel_input         : in    std_logic;
          I_1_RNI3I3E3          : out   std_logic;
          raddr_add1            : in    std_logic;
          HRESETn_c             : in    std_logic;
          HCLK_c                : in    std_logic;
          raddr_rst             : in    std_logic
        );

end RAM_CTRLR_v2;

architecture DEF_ARCH of RAM_CTRLR_v2 is 

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component syncram_2pZ0
    port( alu_sample_10               : out   std_logic;
          alu_sample_0                : out   std_logic;
          alu_sample_1                : out   std_logic;
          reg_sample_in_RNIFA3C       : in    std_logic_vector(15 to 15) := (others => 'U');
          reg_sample_in               : in    std_logic_vector(6 downto 5) := (others => 'U');
          ram_output_1                : out   std_logic;
          ram_output_3                : out   std_logic;
          ram_output_4                : out   std_logic;
          ram_output_5                : out   std_logic;
          ram_output_6                : out   std_logic;
          ram_output_7                : out   std_logic;
          ram_output_8                : out   std_logic;
          ram_output_9                : out   std_logic;
          ram_output_10               : out   std_logic;
          ram_output_11               : out   std_logic;
          ram_output_12               : out   std_logic;
          ram_output_13               : out   std_logic;
          ram_output_14               : out   std_logic;
          ram_output_15               : out   std_logic;
          ram_output_17               : out   std_logic;
          ram_output_0                : out   std_logic;
          ram_output_16               : out   std_logic;
          DIN_REG1                    : out   std_logic_vector(15 to 15);
          counter                     : in    std_logic_vector(7 downto 0) := (others => 'U');
          ram_input                   : in    std_logic_vector(17 downto 0) := (others => 'U');
          I_1_RNI3I3E3                : out   std_logic;
          alu_sel_input               : in    std_logic := 'U';
          HCLK_c                      : in    std_logic := 'U';
          ram_write                   : in    std_logic := 'U';
          ADD_8x8_medium_area_I0_S_0  : in    std_logic := 'U';
          ADD_8x8_medium_area_I24_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I25_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I26_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I27_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I28_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I29_Y_0 : in    std_logic := 'U';
          ADD_8x8_medium_area_I30_Y_0 : in    std_logic := 'U';
          syncram_2pZ0_GND            : in    std_logic := 'U';
          syncram_2pZ0_VCC            : in    std_logic := 'U';
          ram_write_i                 : in    std_logic := 'U'
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_TMP[0]\, \counter[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, \counter[4]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, \counter[2]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, \counter[6]_net_1\, 
        ADD_8x8_medium_area_I20_Y_0, \counter[5]_net_1\, N_5_i, 
        ADD_8x8_medium_area_I20_un1_Y_0, N125_i, 
        ADD_8x8_medium_area_I13_Y_0, \counter[3]_net_1\, 
        ADD_8x8_medium_area_I13_un1_Y_0, 
        ADD_8x8_medium_area_I30_Y_0, \counter[7]_net_1\, N149, 
        ADD_8x8_medium_area_I29_Y_0, N147, 
        ADD_8x8_medium_area_I27_Y_0, N145_i, N135_i, 
        ADD_8x8_medium_area_I24_Y_0, N116, 
        ADD_8x8_medium_area_I25_Y_0, ADD_8x8_medium_area_I28_Y_0, 
        N124, \counter[0]_net_1\, N120, 
        ADD_8x8_medium_area_I0_S_0, ADD_8x8_medium_area_I26_Y_0, 
        N121, \counter_3[7]\, I_34, \counter_3[6]\, I_30, 
        \counter_3[5]\, I_33, \counter_3[4]\, I_28, 
        \counter_3[3]\, I_31, \counter_3[2]\, I_32, 
        \counter_3[1]\, I_27, \counter_3[0]\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

    for all : syncram_2pZ0
	Use entity work.syncram_2pZ0(DEF_ARCH);
begin 


    un1_counter_1_ADD_8x8_medium_area_I20_Y_0 : OA1
      port map(A => \counter[4]_net_1\, B => \counter[5]_net_1\, 
        C => N_5_i, Y => ADD_8x8_medium_area_I20_Y_0);
    
    un1_counter_I_45 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \counter[6]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    un1_counter_I_31 : XOR2
      port map(A => \counter[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_31);
    
    un1_counter_I_36 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    un1_counter_1_ADD_8x8_medium_area_I12_Y : MX2B
      port map(A => N116, B => N_5_i, S => \counter[1]_net_1\, Y
         => N135_i);
    
    un1_counter_1_ADD_8x8_medium_area_I13_Y_0 : OAI1
      port map(A => \counter[2]_net_1\, B => \counter[3]_net_1\, 
        C => N_5_i, Y => ADD_8x8_medium_area_I13_Y_0);
    
    un1_counter_I_44 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \counter[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \counter[2]\ : DFN1C0
      port map(D => \counter_3[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[2]_net_1\);
    
    \counter[7]\ : DFN1C0
      port map(D => \counter_3[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[7]_net_1\);
    
    un1_counter_1_ADD_8x8_medium_area_I29_Y_0 : XNOR3
      port map(A => N_5_i, B => \counter[6]_net_1\, C => N147, Y
         => ADD_8x8_medium_area_I29_Y_0);
    
    un1_counter_I_48 : AND2
      port map(A => \counter[4]_net_1\, B => \counter[5]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    un1_counter_1_ADD_8x8_medium_area_I20_Y : OA1B
      port map(A => N145_i, B => ADD_8x8_medium_area_I20_un1_Y_0, 
        C => ADD_8x8_medium_area_I20_Y_0, Y => N147);
    
    \counter_RNO[0]\ : NOR2A
      port map(A => \DWACT_ADD_CI_0_partial_sum[0]\, B => 
        raddr_rst, Y => \counter_3[0]\);
    
    \counter[6]\ : DFN1C0
      port map(D => \counter_3[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[6]_net_1\);
    
    \counter_RNO[4]\ : NOR2A
      port map(A => I_28, B => raddr_rst, Y => \counter_3[4]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \memRAM.SRAM\ : syncram_2pZ0
      port map(alu_sample_10 => alu_sample_10, alu_sample_0 => 
        alu_sample_0, alu_sample_1 => alu_sample_1, 
        reg_sample_in_RNIFA3C(15) => reg_sample_in_RNIFA3C(15), 
        reg_sample_in(6) => reg_sample_in(6), reg_sample_in(5)
         => reg_sample_in(5), ram_output_1 => ram_output_1, 
        ram_output_3 => ram_output_3, ram_output_4 => 
        ram_output_4, ram_output_5 => ram_output_5, ram_output_6
         => ram_output_6, ram_output_7 => ram_output_7, 
        ram_output_8 => ram_output_8, ram_output_9 => 
        ram_output_9, ram_output_10 => ram_output_10, 
        ram_output_11 => ram_output_11, ram_output_12 => 
        ram_output_12, ram_output_13 => ram_output_13, 
        ram_output_14 => ram_output_14, ram_output_15 => 
        ram_output_15, ram_output_17 => ram_output_17, 
        ram_output_0 => ram_output_0, ram_output_16 => 
        ram_output_16, DIN_REG1(15) => DIN_REG1(15), counter(7)
         => \counter[7]_net_1\, counter(6) => \counter[6]_net_1\, 
        counter(5) => \counter[5]_net_1\, counter(4) => 
        \counter[4]_net_1\, counter(3) => \counter[3]_net_1\, 
        counter(2) => \counter[2]_net_1\, counter(1) => 
        \counter[1]_net_1\, counter(0) => \counter[0]_net_1\, 
        ram_input(17) => ram_input(17), ram_input(16) => 
        ram_input(16), ram_input(15) => ram_input(15), 
        ram_input(14) => ram_input(14), ram_input(13) => 
        ram_input(13), ram_input(12) => ram_input(12), 
        ram_input(11) => ram_input(11), ram_input(10) => 
        ram_input(10), ram_input(9) => ram_input(9), ram_input(8)
         => ram_input(8), ram_input(7) => ram_input(7), 
        ram_input(6) => ram_input(6), ram_input(5) => 
        ram_input(5), ram_input(4) => ram_input(4), ram_input(3)
         => ram_input(3), ram_input(2) => ram_input(2), 
        ram_input(1) => ram_input(1), ram_input(0) => 
        ram_input(0), I_1_RNI3I3E3 => I_1_RNI3I3E3, alu_sel_input
         => alu_sel_input, HCLK_c => HCLK_c, ram_write => 
        ram_write, ADD_8x8_medium_area_I0_S_0 => 
        ADD_8x8_medium_area_I0_S_0, ADD_8x8_medium_area_I24_Y_0
         => ADD_8x8_medium_area_I24_Y_0, 
        ADD_8x8_medium_area_I25_Y_0 => 
        ADD_8x8_medium_area_I25_Y_0, ADD_8x8_medium_area_I26_Y_0
         => ADD_8x8_medium_area_I26_Y_0, 
        ADD_8x8_medium_area_I27_Y_0 => 
        ADD_8x8_medium_area_I27_Y_0, ADD_8x8_medium_area_I28_Y_0
         => ADD_8x8_medium_area_I28_Y_0, 
        ADD_8x8_medium_area_I29_Y_0 => 
        ADD_8x8_medium_area_I29_Y_0, ADD_8x8_medium_area_I30_Y_0
         => ADD_8x8_medium_area_I30_Y_0, syncram_2pZ0_GND => 
        RAM_CTRLR_v2_GND, syncram_2pZ0_VCC => RAM_CTRLR_v2_VCC, 
        ram_write_i => ram_write_i);
    
    un1_counter_1_ADD_8x8_medium_area_I26_Y_0 : AX1E
      port map(A => N120, B => N135_i, C => N121, Y => 
        ADD_8x8_medium_area_I26_Y_0);
    
    \counter_RNO[1]\ : NOR2A
      port map(A => I_27, B => raddr_rst, Y => \counter_3[1]\);
    
    un1_counter_1_ADD_8x8_medium_area_I0_CO1 : OR3B
      port map(A => waddr_previous(0), B => \counter[0]_net_1\, C
         => waddr_previous(1), Y => N116);
    
    \un2_waddr_0_x2[6]\ : XOR2
      port map(A => waddr_previous(1), B => waddr_previous(0), Y
         => N_5_i);
    
    un1_counter_1_ADD_8x8_medium_area_I4_CO1 : OR2B
      port map(A => \counter[4]_net_1\, B => N_5_i, Y => N124);
    
    un1_counter_I_28 : XOR2
      port map(A => \counter[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_28);
    
    un1_counter_1_ADD_8x8_medium_area_I3_S_0 : XOR2
      port map(A => \counter[3]_net_1\, B => N_5_i, Y => N121);
    
    un1_counter_1_ADD_8x8_medium_area_I25_Y_0 : XNOR3
      port map(A => N_5_i, B => \counter[2]_net_1\, C => N135_i, 
        Y => ADD_8x8_medium_area_I25_Y_0);
    
    un1_counter_I_42 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \counter[4]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    un1_counter_1_ADD_8x8_medium_area_I30_Y_0 : XOR3
      port map(A => N_5_i, B => \counter[7]_net_1\, C => N149, Y
         => ADD_8x8_medium_area_I30_Y_0);
    
    un1_counter_I_35 : NOR2B
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \counter[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \counter[4]\ : DFN1C0
      port map(D => \counter_3[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[4]_net_1\);
    
    un1_counter_1_ADD_8x8_medium_area_I20_un1_Y_0 : OR2
      port map(A => \counter[4]_net_1\, B => N125_i, Y => 
        ADD_8x8_medium_area_I20_un1_Y_0);
    
    \counter[5]\ : DFN1C0
      port map(D => \counter_3[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[5]_net_1\);
    
    un1_counter_I_34 : XOR2
      port map(A => \counter[7]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_34);
    
    un1_counter_1_ADD_8x8_medium_area_I21_Y : MX2A
      port map(A => N147, B => N_5_i, S => \counter[6]_net_1\, Y
         => N149);
    
    \counter_RNO[2]\ : NOR2A
      port map(A => I_32, B => raddr_rst, Y => \counter_3[2]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_counter_I_30 : XOR2
      port map(A => \counter[6]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_30);
    
    \counter_RNO[5]\ : NOR2A
      port map(A => I_33, B => raddr_rst, Y => \counter_3[5]\);
    
    \counter_RNO[3]\ : NOR2A
      port map(A => I_31, B => raddr_rst, Y => \counter_3[3]\);
    
    un1_counter_1_ADD_8x8_medium_area_I13_un1_Y_0 : OR2
      port map(A => \counter[2]_net_1\, B => \counter[3]_net_1\, 
        Y => ADD_8x8_medium_area_I13_un1_Y_0);
    
    \counter[1]\ : DFN1C0
      port map(D => \counter_3[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[1]_net_1\);
    
    \counter[3]\ : DFN1C0
      port map(D => \counter_3[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[3]_net_1\);
    
    un1_counter_I_39 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    un1_counter_1_ADD_8x8_medium_area_I0_S_0 : AX1
      port map(A => waddr_previous(1), B => waddr_previous(0), C
         => \counter[0]_net_1\, Y => ADD_8x8_medium_area_I0_S_0);
    
    un1_counter_I_47 : AND2
      port map(A => \counter[2]_net_1\, B => \counter[3]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    un1_counter_I_19 : XOR2
      port map(A => \counter[0]_net_1\, B => raddr_add1, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \counter_RNO[6]\ : NOR2A
      port map(A => I_30, B => raddr_rst, Y => \counter_3[6]\);
    
    un1_counter_I_1 : AND2
      port map(A => \counter[0]_net_1\, B => raddr_add1, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    un1_counter_1_ADD_8x8_medium_area_I5_S_0 : XNOR2
      port map(A => \counter[5]_net_1\, B => N_5_i, Y => N125_i);
    
    un1_counter_1_ADD_8x8_medium_area_I13_Y : OA1
      port map(A => N135_i, B => ADD_8x8_medium_area_I13_un1_Y_0, 
        C => ADD_8x8_medium_area_I13_Y_0, Y => N145_i);
    
    un1_counter_I_33 : XOR2
      port map(A => \counter[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => I_33);
    
    un1_counter_I_32 : XOR2
      port map(A => \counter[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_32);
    
    un1_counter_I_27 : XOR2
      port map(A => \counter[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_27);
    
    un1_counter_1_ADD_8x8_medium_area_I27_Y_0 : XNOR3
      port map(A => N_5_i, B => \counter[4]_net_1\, C => N145_i, 
        Y => ADD_8x8_medium_area_I27_Y_0);
    
    un1_counter_1_ADD_8x8_medium_area_I28_Y_0 : AX1C
      port map(A => N124, B => N145_i, C => N125_i, Y => 
        ADD_8x8_medium_area_I28_Y_0);
    
    un1_counter_1_ADD_8x8_medium_area_I24_Y_0 : XNOR3
      port map(A => N116, B => \counter[1]_net_1\, C => N_5_i, Y
         => ADD_8x8_medium_area_I24_Y_0);
    
    \counter_RNO[7]\ : NOR2A
      port map(A => I_34, B => raddr_rst, Y => \counter_3[7]\);
    
    un1_counter_1_ADD_8x8_medium_area_I2_CO1 : OR2B
      port map(A => \counter[2]_net_1\, B => N_5_i, Y => N120);
    
    \counter[0]\ : DFN1C0
      port map(D => \counter_3[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \counter[0]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity IIR_CEL_CTRLR_v2_DATAFLOW is

    port( alu_ctrl                      : in    std_logic_vector(2 downto 0);
          S                             : out   std_logic_vector(8 to 8);
          S_i_0                         : out   std_logic_vector(33 to 33);
          alu_sel_coeff                 : in    std_logic_vector(4 downto 0);
          alu_sel_coeff_0_2             : in    std_logic;
          alu_sel_coeff_0_0             : in    std_logic;
          waddr_previous                : in    std_logic_vector(1 downto 0);
          sample_0                      : in    std_logic_vector(14 downto 0);
          sample_in_buf                 : in    std_logic_vector(143 downto 129);
          ram_sel_Wdata                 : in    std_logic_vector(1 downto 0);
          sample_out_s_0                : out   std_logic;
          sample_out_s_1                : out   std_logic;
          sample_out_s_3                : out   std_logic;
          sample_out_s_2                : out   std_logic;
          sample_out_s_10               : out   std_logic;
          sample_out_s_15               : out   std_logic;
          sample_out_s_14               : out   std_logic;
          sample_out_s_13               : out   std_logic;
          sample_out_s_12               : out   std_logic;
          sample_out_s_11               : out   std_logic;
          sample_out_s_9                : out   std_logic;
          sample_out_s_8                : out   std_logic;
          sample_out_s_7                : out   std_logic;
          sample_out_s_6                : out   std_logic;
          sample_out_s_5                : out   std_logic;
          sample_out_s_4                : out   std_logic;
          sample_in_s_1                 : in    std_logic_vector(17 to 17);
          in_sel_src                    : in    std_logic_vector(1 downto 0);
          raddr_rst                     : in    std_logic;
          raddr_add1                    : in    std_logic;
          ram_write                     : in    std_logic;
          IIR_CEL_CTRLR_v2_DATAFLOW_GND : in    std_logic;
          IIR_CEL_CTRLR_v2_DATAFLOW_VCC : in    std_logic;
          ram_write_i                   : in    std_logic;
          HRESETn_c                     : in    std_logic;
          HCLK_c                        : in    std_logic;
          sample_val_delay              : in    std_logic;
          alu_sel_input                 : in    std_logic
        );

end IIR_CEL_CTRLR_v2_DATAFLOW;

architecture DEF_ARCH of IIR_CEL_CTRLR_v2_DATAFLOW is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component MUXN_9_5
    port( alu_sel_coeff_0_0 : in    std_logic := 'U';
          alu_sel_coeff_0_2 : in    std_logic := 'U';
          alu_sel_coeff     : in    std_logic_vector(4 downto 0) := (others => 'U');
          S_i_0             : out   std_logic_vector(33 to 33);
          S                 : out   std_logic_vector(8 to 8);
          alu_coef_s        : out   std_logic_vector(8 downto 0)
        );
  end component;

  component ALU
    port( alu_ctrl     : in    std_logic_vector(2 downto 0) := (others => 'U');
          alu_coef_s   : in    std_logic_vector(8 downto 0) := (others => 'U');
          alu_sample   : in    std_logic_vector(17 downto 0) := (others => 'U');
          sample_out_s : out   std_logic_vector(17 downto 0);
          HRESETn_c    : in    std_logic := 'U';
          HCLK_c       : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM_CTRLR_v2
    port( ram_input             : in    std_logic_vector(17 downto 0) := (others => 'U');
          DIN_REG1              : out   std_logic_vector(15 to 15);
          ram_output_16         : out   std_logic;
          ram_output_0          : out   std_logic;
          ram_output_17         : out   std_logic;
          ram_output_15         : out   std_logic;
          ram_output_14         : out   std_logic;
          ram_output_13         : out   std_logic;
          ram_output_12         : out   std_logic;
          ram_output_11         : out   std_logic;
          ram_output_10         : out   std_logic;
          ram_output_9          : out   std_logic;
          ram_output_8          : out   std_logic;
          ram_output_7          : out   std_logic;
          ram_output_6          : out   std_logic;
          ram_output_5          : out   std_logic;
          ram_output_4          : out   std_logic;
          ram_output_3          : out   std_logic;
          ram_output_1          : out   std_logic;
          reg_sample_in         : in    std_logic_vector(6 downto 5) := (others => 'U');
          reg_sample_in_RNIFA3C : in    std_logic_vector(15 to 15) := (others => 'U');
          alu_sample_1          : out   std_logic;
          alu_sample_0          : out   std_logic;
          alu_sample_10         : out   std_logic;
          waddr_previous        : in    std_logic_vector(1 downto 0) := (others => 'U');
          ram_write_i           : in    std_logic := 'U';
          RAM_CTRLR_v2_VCC      : in    std_logic := 'U';
          RAM_CTRLR_v2_GND      : in    std_logic := 'U';
          ram_write             : in    std_logic := 'U';
          alu_sel_input         : in    std_logic := 'U';
          I_1_RNI3I3E3          : out   std_logic;
          raddr_add1            : in    std_logic := 'U';
          HRESETn_c             : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U';
          raddr_rst             : in    std_logic := 'U'
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \reg_sample_in_RNIFA3C[15]_net_1\, 
        \reg_sample_in[15]_net_1\, \DIN_REG1[15]\, 
        \reg_sample_in6\, N_318, \ram_output[4]\, 
        \sample_in_s_27[4]\, N_319, \ram_output[5]\, 
        \sample_in_s_25[5]\, N_320, \ram_output[6]\, 
        \sample_in_s_23[6]\, N_321, \ram_output[7]\, 
        \sample_in_s_21[7]\, N_322, \ram_output[8]\, 
        \sample_in_s_19[8]\, N_323, \ram_output[9]\, 
        \sample_in_s_17[9]\, N_324, \ram_output[10]\, 
        \sample_in_s_15[10]\, N_325, \ram_output[11]\, 
        \sample_in_s_13[11]\, N_326, \ram_output[12]\, 
        \sample_in_s_11[12]\, N_327, \ram_output[13]\, 
        \sample_in_s_9[13]\, N_328, \ram_output[14]\, 
        \sample_in_s_7[14]\, N_329, \ram_output[15]\, N_331, 
        \ram_output[17]\, \reg_sample_in_5[4]\, 
        reg_sample_in_5_sn_N_2_i, \reg_sample_in_5[5]\, 
        \reg_sample_in_5[6]\, \reg_sample_in_5[7]\, 
        \reg_sample_in_5[8]\, \reg_sample_in_5[9]\, 
        \reg_sample_in_5[11]\, \reg_sample_in_5[12]\, 
        \reg_sample_in_5[13]\, \reg_sample_in_5[14]\, 
        \reg_sample_in_5[15]\, \reg_sample_in_5[17]\, 
        \sample_out_s[17]\, N_358, \reg_sample_in[4]_net_1\, 
        \sample_out_s[4]\, N_359, \reg_sample_in[5]_net_1\, 
        \sample_out_s[5]\, N_360, \reg_sample_in[6]_net_1\, 
        \sample_out_s[6]\, N_361, \reg_sample_in[7]_net_1\, 
        \sample_out_s[7]\, N_362, \reg_sample_in[8]_net_1\, 
        \sample_out_s[8]\, N_363, \reg_sample_in[9]_net_1\, 
        \sample_out_s[9]\, N_364, \reg_sample_in[10]_net_1\, 
        N_365, \reg_sample_in[11]_net_1\, \sample_out_s[11]\, 
        N_366, \reg_sample_in[12]_net_1\, \sample_out_s[12]\, 
        N_367, \reg_sample_in[13]_net_1\, \sample_out_s[13]\, 
        N_368, \reg_sample_in[14]_net_1\, \sample_out_s[14]\, 
        N_369, \sample_out_s[15]\, N_371, 
        \reg_sample_in[17]_net_1\, \ram_input[4]\, \ram_input[5]\, 
        \ram_input[6]\, \ram_input[7]\, \ram_input[8]\, 
        \ram_input[9]\, \ram_input[10]\, \ram_input[11]\, 
        \ram_input[12]\, \ram_input[13]\, \ram_input[14]\, 
        \ram_input[15]\, \ram_input[17]\, \alu_sample[1]\, 
        \reg_sample_in[1]_net_1\, \ram_output[1]\, 
        \alu_sample[2]\, \reg_sample_in[2]_net_1\, I_1_RNI3I3E3, 
        \alu_sample[3]\, \reg_sample_in[3]_net_1\, 
        \ram_output[3]\, \alu_sample[4]\, \alu_sample[7]\, 
        \alu_sample[8]\, \alu_sample[9]\, \alu_sample[11]\, 
        \alu_sample[12]\, \alu_sample[13]\, \alu_sample[14]\, 
        \alu_sample[17]\, N_316, \sample_in_s_31[2]\, N_317, 
        \sample_in_s_29[3]\, \reg_sample_in_5[2]\, 
        \reg_sample_in_5[3]\, N_356, \sample_out_s[2]\, N_357, 
        \sample_out_s[3]\, \ram_input[2]\, \ram_input[3]\, N_315, 
        \sample_in_s_33[1]\, \reg_sample_in_5[1]\, N_355, 
        \sample_out_s[1]\, \ram_input[1]\, \alu_sample[10]\, 
        \reg_sample_in_5[10]\, \sample_out_s[10]\, 
        \sample_in_s_35[0]\, \ram_input[0]\, N_354, 
        \ram_output[0]\, \reg_sample_in[0]_net_1\, 
        \reg_sample_in_5[0]\, \sample_out_s[0]\, N_314, 
        \alu_sample[0]\, \alu_sample[16]\, 
        \reg_sample_in[16]_net_1\, \ram_output[16]\, 
        \ram_input[16]\, N_370, \sample_out_s[16]\, 
        \reg_sample_in_5[16]\, N_330, \alu_sample[6]\, 
        \alu_sample[5]\, \alu_sample[15]\, \alu_coef_s[0]\, 
        \alu_coef_s[1]\, \alu_coef_s[2]\, \alu_coef_s[3]\, 
        \alu_coef_s[4]\, \alu_coef_s[5]\, \alu_coef_s[6]\, 
        \alu_coef_s[7]\, \alu_coef_s[8]\, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

    for all : MUXN_9_5
	Use entity work.MUXN_9_5(DEF_ARCH);
    for all : ALU
	Use entity work.ALU(DEF_ARCH);
    for all : RAM_CTRLR_v2
	Use entity work.RAM_CTRLR_v2(DEF_ARCH);
begin 

    sample_out_s_0 <= \sample_out_s[0]\;
    sample_out_s_1 <= \sample_out_s[1]\;
    sample_out_s_3 <= \sample_out_s[3]\;
    sample_out_s_2 <= \sample_out_s[2]\;
    sample_out_s_10 <= \sample_out_s[10]\;
    sample_out_s_15 <= \sample_out_s[15]\;
    sample_out_s_14 <= \sample_out_s[14]\;
    sample_out_s_13 <= \sample_out_s[13]\;
    sample_out_s_12 <= \sample_out_s[12]\;
    sample_out_s_11 <= \sample_out_s[11]\;
    sample_out_s_9 <= \sample_out_s[9]\;
    sample_out_s_8 <= \sample_out_s[8]\;
    sample_out_s_7 <= \sample_out_s[7]\;
    sample_out_s_6 <= \sample_out_s[6]\;
    sample_out_s_5 <= \sample_out_s[5]\;
    sample_out_s_4 <= \sample_out_s[4]\;

    \reg_sample_in_RNO_1[10]\ : MX2
      port map(A => sample_in_buf(133), B => sample_0(10), S => 
        sample_val_delay, Y => \sample_in_s_15[10]\);
    
    \reg_sample_in_RNO[2]\ : MX2
      port map(A => \sample_out_s[2]\, B => N_316, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[2]\);
    
    \reg_sample_in_RNIO8MA4[8]\ : MX2
      port map(A => N_362, B => \ram_output[8]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[8]\);
    
    \reg_sample_in_RNO_1[1]\ : MX2
      port map(A => sample_in_buf(142), B => sample_0(1), S => 
        sample_val_delay, Y => \sample_in_s_33[1]\);
    
    \reg_sample_in_RNIUJBJ[12]\ : MX2
      port map(A => \reg_sample_in[12]_net_1\, B => 
        \sample_out_s[12]\, S => ram_sel_Wdata(0), Y => N_366);
    
    \reg_sample_in_RNIJLRL3[11]\ : MX2
      port map(A => \reg_sample_in[11]_net_1\, B => 
        \ram_output[11]\, S => alu_sel_input, Y => 
        \alu_sample[11]\);
    
    \reg_sample_in_RNO_0[7]\ : MX2
      port map(A => \ram_output[7]\, B => \sample_in_s_21[7]\, S
         => in_sel_src(0), Y => N_321);
    
    \reg_sample_in_RNIPLRL3[14]\ : MX2
      port map(A => \reg_sample_in[14]_net_1\, B => 
        \ram_output[14]\, S => alu_sel_input, Y => 
        \alu_sample[14]\);
    
    \reg_sample_in_RNII1984[2]\ : MX2
      port map(A => N_356, B => I_1_RNI3I3E3, S => 
        ram_sel_Wdata(1), Y => \ram_input[2]\);
    
    \reg_sample_in[5]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[5]_net_1\);
    
    \reg_sample_in_RNI0HPO[5]\ : MX2C
      port map(A => \reg_sample_in[5]_net_1\, B => 
        \sample_out_s[5]\, S => ram_sel_Wdata(0), Y => N_359);
    
    \reg_sample_in_RNISOMA4[9]\ : MX2
      port map(A => N_363, B => \ram_output[9]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[9]\);
    
    \reg_sample_in_RNI1U5Q3[0]\ : MX2
      port map(A => \reg_sample_in[0]_net_1\, B => 
        \ram_output[0]\, S => alu_sel_input, Y => \alu_sample[0]\);
    
    \reg_sample_in_RNIJ68Q3[9]\ : MX2
      port map(A => \reg_sample_in[9]_net_1\, B => 
        \ram_output[9]\, S => alu_sel_input, Y => \alu_sample[9]\);
    
    \reg_sample_in_RNI4OJA4[3]\ : MX2
      port map(A => N_357, B => \ram_output[3]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[3]\);
    
    \reg_sample_in_RNO_0[0]\ : MX2
      port map(A => \ram_output[0]\, B => \sample_in_s_35[0]\, S
         => in_sel_src(0), Y => N_314);
    
    \reg_sample_in_RNO_0[1]\ : MX2
      port map(A => \ram_output[1]\, B => \sample_in_s_33[1]\, S
         => in_sel_src(0), Y => N_315);
    
    \reg_sample_in_RNI3TPO[6]\ : MX2C
      port map(A => \reg_sample_in[6]_net_1\, B => 
        \sample_out_s[6]\, S => ram_sel_Wdata(0), Y => N_360);
    
    \reg_sample_in_RNO_0[2]\ : MX2
      port map(A => I_1_RNI3I3E3, B => \sample_in_s_31[2]\, S => 
        in_sel_src(0), Y => N_316);
    
    \reg_sample_in_RNIT4PO[4]\ : MX2
      port map(A => \reg_sample_in[4]_net_1\, B => 
        \sample_out_s[4]\, S => ram_sel_Wdata(0), Y => N_358);
    
    \reg_sample_in_RNO[11]\ : MX2
      port map(A => \sample_out_s[11]\, B => N_325, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[11]\);
    
    \reg_sample_in_RNO_1[2]\ : MX2
      port map(A => sample_in_buf(141), B => sample_0(2), S => 
        sample_val_delay, Y => \sample_in_s_31[2]\);
    
    \reg_sample_in_RNO_0[11]\ : MX2
      port map(A => \ram_output[11]\, B => \sample_in_s_13[11]\, 
        S => in_sel_src(0), Y => N_325);
    
    \reg_sample_in_RNIU7964[15]\ : MX2
      port map(A => N_369, B => \ram_output[15]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[15]\);
    
    reg_sample_in6 : NOR2
      port map(A => in_sel_src(1), B => in_sel_src(0), Y => 
        \reg_sample_in6\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \reg_sample_in_RNO[13]\ : MX2
      port map(A => \sample_out_s[13]\, B => N_327, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[13]\);
    
    \reg_sample_in[3]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[3]_net_1\);
    
    \reg_sample_in_RNO_1[9]\ : MX2
      port map(A => sample_in_buf(134), B => sample_0(9), S => 
        sample_val_delay, Y => \sample_in_s_17[9]\);
    
    \reg_sample_in_RNO[4]\ : MX2
      port map(A => \sample_out_s[4]\, B => N_318, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[4]\);
    
    \reg_sample_in[7]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[7]_net_1\);
    
    \reg_sample_in[14]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[14]_net_1\);
    
    \reg_sample_in_RNILLRL3[12]\ : MX2
      port map(A => \reg_sample_in[12]_net_1\, B => 
        \ram_output[12]\, S => alu_sel_input, Y => 
        \alu_sample[12]\);
    
    \reg_sample_in_RNIEP884[1]\ : MX2
      port map(A => N_355, B => \ram_output[1]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[1]\);
    
    \reg_sample_in_RNO[3]\ : MX2
      port map(A => \sample_out_s[3]\, B => N_317, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[3]\);
    
    \reg_sample_in_RNI5E6Q3[2]\ : MX2
      port map(A => \reg_sample_in[2]_net_1\, B => I_1_RNI3I3E3, 
        S => alu_sel_input, Y => \alu_sample[2]\);
    
    \reg_sample_in_RNO_1[11]\ : MX2
      port map(A => sample_in_buf(132), B => sample_0(11), S => 
        sample_val_delay, Y => \sample_in_s_13[11]\);
    
    \reg_sample_in_RNO[1]\ : MX2
      port map(A => \sample_out_s[1]\, B => N_315, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[1]\);
    
    \reg_sample_in_RNI9U6Q3[4]\ : MX2
      port map(A => \reg_sample_in[4]_net_1\, B => 
        \ram_output[4]\, S => alu_sel_input, Y => \alu_sample[4]\);
    
    \reg_sample_in[9]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[9]_net_1\);
    
    \reg_sample_in_RNO_0[15]\ : MX2
      port map(A => \ram_output[15]\, B => sample_in_s_1(17), S
         => in_sel_src(0), Y => N_329);
    
    \reg_sample_in_RNO[8]\ : MX2
      port map(A => \sample_out_s[8]\, B => N_322, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[8]\);
    
    \reg_sample_in_RNO[12]\ : MX2
      port map(A => \sample_out_s[12]\, B => N_326, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[12]\);
    
    \reg_sample_in_RNI6O964[17]\ : MX2
      port map(A => N_371, B => \ram_output[17]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[17]\);
    
    \reg_sample_in_RNIFB9J[13]\ : MX2
      port map(A => \reg_sample_in[13]_net_1\, B => 
        \sample_out_s[13]\, S => ram_sel_Wdata(0), Y => N_367);
    
    \reg_sample_in_RNIRBBJ[11]\ : MX2
      port map(A => \reg_sample_in[11]_net_1\, B => 
        \sample_out_s[11]\, S => ram_sel_Wdata(0), Y => N_365);
    
    \reg_sample_in_RNIQOOO[3]\ : MX2
      port map(A => \reg_sample_in[3]_net_1\, B => 
        \sample_out_s[3]\, S => ram_sel_Wdata(0), Y => N_357);
    
    \reg_sample_in_RNIFA3C[15]\ : MX2
      port map(A => \reg_sample_in[15]_net_1\, B => 
        \DIN_REG1[15]\, S => alu_sel_input, Y => 
        \reg_sample_in_RNIFA3C[15]_net_1\);
    
    \reg_sample_in_RNI0OA64[11]\ : MX2
      port map(A => N_365, B => \ram_output[11]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[11]\);
    
    \reg_sample_in_RNO_0[16]\ : MX2
      port map(A => \ram_output[16]\, B => sample_in_s_1(17), S
         => in_sel_src(0), Y => N_330);
    
    \reg_sample_in_RNIIJ9J[14]\ : MX2
      port map(A => \reg_sample_in[14]_net_1\, B => 
        \sample_out_s[14]\, S => ram_sel_Wdata(0), Y => N_368);
    
    \reg_sample_in[16]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[16]_net_1\);
    
    \reg_sample_in_RNO_1[5]\ : MX2C
      port map(A => sample_in_buf(138), B => sample_0(5), S => 
        sample_val_delay, Y => \sample_in_s_25[5]\);
    
    \reg_sample_in_RNIVLRL3[17]\ : MX2
      port map(A => \reg_sample_in[17]_net_1\, B => 
        \ram_output[17]\, S => alu_sel_input, Y => 
        \alu_sample[17]\);
    
    \reg_sample_in_RNIFM7Q3[7]\ : MX2
      port map(A => \reg_sample_in[7]_net_1\, B => 
        \ram_output[7]\, S => alu_sel_input, Y => \alu_sample[7]\);
    
    Coeff_Mux : MUXN_9_5
      port map(alu_sel_coeff_0_0 => alu_sel_coeff_0_0, 
        alu_sel_coeff_0_2 => alu_sel_coeff_0_2, alu_sel_coeff(4)
         => alu_sel_coeff(4), alu_sel_coeff(3) => 
        alu_sel_coeff(3), alu_sel_coeff(2) => alu_sel_coeff(2), 
        alu_sel_coeff(1) => alu_sel_coeff(1), alu_sel_coeff(0)
         => alu_sel_coeff(0), S_i_0(33) => S_i_0(33), S(8) => 
        S(8), alu_coef_s(8) => \alu_coef_s[8]\, alu_coef_s(7) => 
        \alu_coef_s[7]\, alu_coef_s(6) => \alu_coef_s[6]\, 
        alu_coef_s(5) => \alu_coef_s[5]\, alu_coef_s(4) => 
        \alu_coef_s[4]\, alu_coef_s(3) => \alu_coef_s[3]\, 
        alu_coef_s(2) => \alu_coef_s[2]\, alu_coef_s(1) => 
        \alu_coef_s[1]\, alu_coef_s(0) => \alu_coef_s[0]\);
    
    ALU_1 : ALU
      port map(alu_ctrl(2) => alu_ctrl(2), alu_ctrl(1) => 
        alu_ctrl(1), alu_ctrl(0) => alu_ctrl(0), alu_coef_s(8)
         => \alu_coef_s[8]\, alu_coef_s(7) => \alu_coef_s[7]\, 
        alu_coef_s(6) => \alu_coef_s[6]\, alu_coef_s(5) => 
        \alu_coef_s[5]\, alu_coef_s(4) => \alu_coef_s[4]\, 
        alu_coef_s(3) => \alu_coef_s[3]\, alu_coef_s(2) => 
        \alu_coef_s[2]\, alu_coef_s(1) => \alu_coef_s[1]\, 
        alu_coef_s(0) => \alu_coef_s[0]\, alu_sample(17) => 
        \alu_sample[17]\, alu_sample(16) => \alu_sample[16]\, 
        alu_sample(15) => \alu_sample[15]\, alu_sample(14) => 
        \alu_sample[14]\, alu_sample(13) => \alu_sample[13]\, 
        alu_sample(12) => \alu_sample[12]\, alu_sample(11) => 
        \alu_sample[11]\, alu_sample(10) => \alu_sample[10]\, 
        alu_sample(9) => \alu_sample[9]\, alu_sample(8) => 
        \alu_sample[8]\, alu_sample(7) => \alu_sample[7]\, 
        alu_sample(6) => \alu_sample[6]\, alu_sample(5) => 
        \alu_sample[5]\, alu_sample(4) => \alu_sample[4]\, 
        alu_sample(3) => \alu_sample[3]\, alu_sample(2) => 
        \alu_sample[2]\, alu_sample(1) => \alu_sample[1]\, 
        alu_sample(0) => \alu_sample[0]\, sample_out_s(17) => 
        \sample_out_s[17]\, sample_out_s(16) => 
        \sample_out_s[16]\, sample_out_s(15) => 
        \sample_out_s[15]\, sample_out_s(14) => 
        \sample_out_s[14]\, sample_out_s(13) => 
        \sample_out_s[13]\, sample_out_s(12) => 
        \sample_out_s[12]\, sample_out_s(11) => 
        \sample_out_s[11]\, sample_out_s(10) => 
        \sample_out_s[10]\, sample_out_s(9) => \sample_out_s[9]\, 
        sample_out_s(8) => \sample_out_s[8]\, sample_out_s(7) => 
        \sample_out_s[7]\, sample_out_s(6) => \sample_out_s[6]\, 
        sample_out_s(5) => \sample_out_s[5]\, sample_out_s(4) => 
        \sample_out_s[4]\, sample_out_s(3) => \sample_out_s[3]\, 
        sample_out_s(2) => \sample_out_s[2]\, sample_out_s(1) => 
        \sample_out_s[1]\, sample_out_s(0) => \sample_out_s[0]\, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c);
    
    \reg_sample_in_RNI7M6Q3[3]\ : MX2
      port map(A => \reg_sample_in[3]_net_1\, B => 
        \ram_output[3]\, S => alu_sel_input, Y => \alu_sample[3]\);
    
    \reg_sample_in[8]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[8]_net_1\);
    
    \reg_sample_in[13]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[13]_net_1\);
    
    \reg_sample_in[12]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[12]_net_1\);
    
    \reg_sample_in_RNISFA64[10]\ : MX2
      port map(A => N_364, B => \ram_output[10]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[10]\);
    
    \reg_sample_in_RNIHLRL3[10]\ : MX2
      port map(A => \reg_sample_in[10]_net_1\, B => 
        \ram_output[10]\, S => alu_sel_input, Y => 
        \alu_sample[10]\);
    
    \reg_sample_in_RNI88KA4[4]\ : MX2
      port map(A => N_358, B => \ram_output[4]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[4]\);
    
    \reg_sample_in_RNI62EM[1]\ : MX2
      port map(A => \reg_sample_in[1]_net_1\, B => 
        \sample_out_s[1]\, S => ram_sel_Wdata(0), Y => N_355);
    
    \reg_sample_in[10]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[10]_net_1\);
    
    \reg_sample_in[6]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[6]_net_1\);
    
    \reg_sample_in[1]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[1]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \reg_sample_in_RNO[10]\ : MX2
      port map(A => \sample_out_s[10]\, B => N_324, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[10]\);
    
    \reg_sample_in_RNIC1RO[9]\ : MX2
      port map(A => \reg_sample_in[9]_net_1\, B => 
        \sample_out_s[9]\, S => ram_sel_Wdata(0), Y => N_363);
    
    \reg_sample_in_RNIQV864[14]\ : MX2
      port map(A => N_368, B => \ram_output[14]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[14]\);
    
    \reg_sample_in_RNIO3AJ[16]\ : MX2
      port map(A => \reg_sample_in[16]_net_1\, B => 
        \sample_out_s[16]\, S => ram_sel_Wdata(0), Y => N_370);
    
    \reg_sample_in_RNO_0[5]\ : MX2C
      port map(A => \ram_output[5]\, B => \sample_in_s_25[5]\, S
         => in_sel_src(0), Y => N_319);
    
    \reg_sample_in_RNIAH884[0]\ : MX2
      port map(A => N_354, B => \ram_output[0]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[0]\);
    
    \reg_sample_in[2]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[2]_net_1\);
    
    \reg_sample_in_RNO_1[4]\ : MX2
      port map(A => sample_in_buf(139), B => sample_0(4), S => 
        sample_val_delay, Y => \sample_in_s_27[4]\);
    
    \reg_sample_in_RNI40B64[12]\ : MX2
      port map(A => N_366, B => \ram_output[12]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[12]\);
    
    \reg_sample_in_RNIO3BJ[10]\ : MX2
      port map(A => \reg_sample_in[10]_net_1\, B => 
        \sample_out_s[10]\, S => ram_sel_Wdata(0), Y => N_364);
    
    \reg_sample_in[17]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[17]_net_1\);
    
    \reg_sample_in_RNO[7]\ : MX2
      port map(A => \sample_out_s[7]\, B => N_321, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[7]\);
    
    \reg_sample_in_RNO[16]\ : MX2
      port map(A => \sample_out_s[16]\, B => N_330, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[16]\);
    
    \reg_sample_in_RNI9LQO[8]\ : MX2
      port map(A => \reg_sample_in[8]_net_1\, B => 
        \sample_out_s[8]\, S => ram_sel_Wdata(0), Y => N_362);
    
    \reg_sample_in[4]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[4]_net_1\);
    
    \reg_sample_in_RNO_1[7]\ : MX2
      port map(A => sample_in_buf(136), B => sample_0(7), S => 
        sample_val_delay, Y => \sample_in_s_21[7]\);
    
    \reg_sample_in_RNO_1[3]\ : MX2
      port map(A => sample_in_buf(140), B => sample_0(3), S => 
        sample_val_delay, Y => \sample_in_s_29[3]\);
    
    \reg_sample_in_RNO_0[12]\ : MX2
      port map(A => \ram_output[12]\, B => \sample_in_s_11[12]\, 
        S => in_sel_src(0), Y => N_326);
    
    \reg_sample_in_RNO[6]\ : MX2
      port map(A => \sample_out_s[6]\, B => N_320, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[6]\);
    
    \reg_sample_in[15]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[15]_net_1\);
    
    \reg_sample_in_RNO_0[4]\ : MX2
      port map(A => \ram_output[4]\, B => \sample_in_s_27[4]\, S
         => in_sel_src(0), Y => N_318);
    
    \reg_sample_in_RNO_0[3]\ : MX2
      port map(A => \ram_output[3]\, B => \sample_in_s_29[3]\, S
         => in_sel_src(0), Y => N_317);
    
    \reg_sample_in_RNO_0[17]\ : MX2
      port map(A => \ram_output[17]\, B => sample_in_s_1(17), S
         => in_sel_src(0), Y => N_331);
    
    \reg_sample_in_RNO[17]\ : MX2
      port map(A => \sample_out_s[17]\, B => N_331, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[17]\);
    
    \reg_sample_in_RNO[14]\ : MX2
      port map(A => \sample_out_s[14]\, B => N_328, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[14]\);
    
    \reg_sample_in_RNIRBAJ[17]\ : MX2
      port map(A => \reg_sample_in[17]_net_1\, B => 
        \sample_out_s[17]\, S => ram_sel_Wdata(0), Y => N_371);
    
    \reg_sample_in_RNO_1[8]\ : MX2
      port map(A => sample_in_buf(135), B => sample_0(8), S => 
        sample_val_delay, Y => \sample_in_s_19[8]\);
    
    \reg_sample_in_RNI3UDM[0]\ : MX2
      port map(A => \reg_sample_in[0]_net_1\, B => 
        \sample_out_s[0]\, S => ram_sel_Wdata(0), Y => N_354);
    
    \reg_sample_in[11]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[11]_net_1\);
    
    \reg_sample_in_RNO[5]\ : MX2
      port map(A => \sample_out_s[5]\, B => N_319, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[5]\);
    
    \reg_sample_in_RNO_0[9]\ : MX2
      port map(A => \ram_output[9]\, B => \sample_in_s_17[9]\, S
         => in_sel_src(0), Y => N_323);
    
    \reg_sample_in_RNO[9]\ : MX2
      port map(A => \sample_out_s[9]\, B => N_323, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[9]\);
    
    RAM_CTRLR_v2_1 : RAM_CTRLR_v2
      port map(ram_input(17) => \ram_input[17]\, ram_input(16)
         => \ram_input[16]\, ram_input(15) => \ram_input[15]\, 
        ram_input(14) => \ram_input[14]\, ram_input(13) => 
        \ram_input[13]\, ram_input(12) => \ram_input[12]\, 
        ram_input(11) => \ram_input[11]\, ram_input(10) => 
        \ram_input[10]\, ram_input(9) => \ram_input[9]\, 
        ram_input(8) => \ram_input[8]\, ram_input(7) => 
        \ram_input[7]\, ram_input(6) => \ram_input[6]\, 
        ram_input(5) => \ram_input[5]\, ram_input(4) => 
        \ram_input[4]\, ram_input(3) => \ram_input[3]\, 
        ram_input(2) => \ram_input[2]\, ram_input(1) => 
        \ram_input[1]\, ram_input(0) => \ram_input[0]\, 
        DIN_REG1(15) => \DIN_REG1[15]\, ram_output_16 => 
        \ram_output[16]\, ram_output_0 => \ram_output[0]\, 
        ram_output_17 => \ram_output[17]\, ram_output_15 => 
        \ram_output[15]\, ram_output_14 => \ram_output[14]\, 
        ram_output_13 => \ram_output[13]\, ram_output_12 => 
        \ram_output[12]\, ram_output_11 => \ram_output[11]\, 
        ram_output_10 => \ram_output[10]\, ram_output_9 => 
        \ram_output[9]\, ram_output_8 => \ram_output[8]\, 
        ram_output_7 => \ram_output[7]\, ram_output_6 => 
        \ram_output[6]\, ram_output_5 => \ram_output[5]\, 
        ram_output_4 => \ram_output[4]\, ram_output_3 => 
        \ram_output[3]\, ram_output_1 => \ram_output[1]\, 
        reg_sample_in(6) => \reg_sample_in[6]_net_1\, 
        reg_sample_in(5) => \reg_sample_in[5]_net_1\, 
        reg_sample_in_RNIFA3C(15) => 
        \reg_sample_in_RNIFA3C[15]_net_1\, alu_sample_1 => 
        \alu_sample[6]\, alu_sample_0 => \alu_sample[5]\, 
        alu_sample_10 => \alu_sample[15]\, waddr_previous(1) => 
        waddr_previous(1), waddr_previous(0) => waddr_previous(0), 
        ram_write_i => ram_write_i, RAM_CTRLR_v2_VCC => 
        IIR_CEL_CTRLR_v2_DATAFLOW_VCC, RAM_CTRLR_v2_GND => 
        IIR_CEL_CTRLR_v2_DATAFLOW_GND, ram_write => ram_write, 
        alu_sel_input => alu_sel_input, I_1_RNI3I3E3 => 
        I_1_RNI3I3E3, raddr_add1 => raddr_add1, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, raddr_rst => raddr_rst);
    
    reg_sample_in_5_sn_m1 : OR2B
      port map(A => in_sel_src(1), B => in_sel_src(0), Y => 
        reg_sample_in_5_sn_N_2_i);
    
    \reg_sample_in_RNO[15]\ : MX2
      port map(A => \sample_out_s[15]\, B => N_329, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[15]\);
    
    \reg_sample_in_RNO_0[14]\ : MX2
      port map(A => \ram_output[14]\, B => \sample_in_s_7[14]\, S
         => in_sel_src(0), Y => N_328);
    
    \reg_sample_in_RNI96EM[2]\ : MX2
      port map(A => \reg_sample_in[2]_net_1\, B => 
        \sample_out_s[2]\, S => ram_sel_Wdata(0), Y => N_356);
    
    \reg_sample_in_RNO_1[12]\ : MX2
      port map(A => sample_in_buf(131), B => sample_0(12), S => 
        sample_val_delay, Y => \sample_in_s_11[12]\);
    
    \reg_sample_in_RNI366Q3[1]\ : MX2
      port map(A => \reg_sample_in[1]_net_1\, B => 
        \ram_output[1]\, S => alu_sel_input, Y => \alu_sample[1]\);
    
    \reg_sample_in_RNI69QO[7]\ : MX2
      port map(A => \reg_sample_in[7]_net_1\, B => 
        \sample_out_s[7]\, S => ram_sel_Wdata(0), Y => N_361);
    
    \reg_sample_in_RNIG8LA4[6]\ : MX2C
      port map(A => N_360, B => \ram_output[6]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[6]\);
    
    \reg_sample_in_RNO_0[8]\ : MX2
      port map(A => \ram_output[8]\, B => \sample_in_s_19[8]\, S
         => in_sel_src(0), Y => N_322);
    
    \reg_sample_in_RNO_0[13]\ : MX2
      port map(A => \ram_output[13]\, B => \sample_in_s_9[13]\, S
         => in_sel_src(0), Y => N_327);
    
    \reg_sample_in_RNO[0]\ : MX2
      port map(A => \sample_out_s[0]\, B => N_314, S => 
        reg_sample_in_5_sn_N_2_i, Y => \reg_sample_in_5[0]\);
    
    \reg_sample_in_RNITLRL3[16]\ : MX2
      port map(A => \reg_sample_in[16]_net_1\, B => 
        \ram_output[16]\, S => alu_sel_input, Y => 
        \alu_sample[16]\);
    
    \reg_sample_in_RNILR9J[15]\ : MX2
      port map(A => \reg_sample_in[15]_net_1\, B => 
        \sample_out_s[15]\, S => ram_sel_Wdata(0), Y => N_369);
    
    \reg_sample_in[0]\ : DFN1E0C0
      port map(D => \reg_sample_in_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \reg_sample_in6\, Q => 
        \reg_sample_in[0]_net_1\);
    
    \reg_sample_in_RNO_0[10]\ : MX2
      port map(A => \ram_output[10]\, B => \sample_in_s_15[10]\, 
        S => in_sel_src(0), Y => N_324);
    
    \reg_sample_in_RNIKOLA4[7]\ : MX2
      port map(A => N_361, B => \ram_output[7]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[7]\);
    
    \reg_sample_in_RNI2G964[16]\ : MX2
      port map(A => N_370, B => \ram_output[16]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[16]\);
    
    \reg_sample_in_RNINLRL3[13]\ : MX2
      port map(A => \reg_sample_in[13]_net_1\, B => 
        \ram_output[13]\, S => alu_sel_input, Y => 
        \alu_sample[13]\);
    
    \reg_sample_in_RNO_1[14]\ : MX2
      port map(A => sample_in_buf(129), B => sample_0(14), S => 
        sample_val_delay, Y => \sample_in_s_7[14]\);
    
    \reg_sample_in_RNO_1[6]\ : MX2C
      port map(A => sample_in_buf(137), B => sample_0(6), S => 
        sample_val_delay, Y => \sample_in_s_23[6]\);
    
    \reg_sample_in_RNIHU7Q3[8]\ : MX2
      port map(A => \reg_sample_in[8]_net_1\, B => 
        \ram_output[8]\, S => alu_sel_input, Y => \alu_sample[8]\);
    
    \reg_sample_in_RNO_0[6]\ : MX2C
      port map(A => \ram_output[6]\, B => \sample_in_s_23[6]\, S
         => in_sel_src(0), Y => N_320);
    
    \reg_sample_in_RNO_1[13]\ : MX2
      port map(A => sample_in_buf(130), B => sample_0(13), S => 
        sample_val_delay, Y => \sample_in_s_9[13]\);
    
    \reg_sample_in_RNO_1[0]\ : MX2
      port map(A => sample_in_buf(143), B => sample_0(0), S => 
        sample_val_delay, Y => \sample_in_s_35[0]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \reg_sample_in_RNIMN864[13]\ : MX2
      port map(A => N_367, B => \ram_output[13]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[13]\);
    
    \reg_sample_in_RNICOKA4[5]\ : MX2C
      port map(A => N_359, B => \ram_output[5]\, S => 
        ram_sel_Wdata(1), Y => \ram_input[5]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity IIR_CEL_CTRLR_v2_CONTROL is

    port( alu_ctrl             : out   std_logic_vector(2 downto 0);
          ram_sel_Wdata        : out   std_logic_vector(1 downto 0);
          waddr_previous       : out   std_logic_vector(1 downto 0);
          in_sel_src           : out   std_logic_vector(1 downto 0);
          S_i_0                : in    std_logic_vector(33 to 33);
          S                    : in    std_logic_vector(8 to 8);
          alu_sel_coeff        : out   std_logic_vector(4 downto 0);
          alu_sel_coeff_0_2    : out   std_logic;
          alu_sel_coeff_0_0    : out   std_logic;
          sample_out_rot_s     : out   std_logic;
          sample_out_val_s     : out   std_logic;
          raddr_rst            : out   std_logic;
          alu_sel_input        : out   std_logic;
          raddr_add1           : out   std_logic;
          sample_val_delay     : in    std_logic;
          ram_write            : out   std_logic;
          ram_write_i          : out   std_logic;
          un1_sample_in_rotate : out   std_logic;
          sample_out_rot_s_0   : out   std_logic;
          sample_out_rot_s_1   : out   std_logic;
          sample_out_rot_s_2   : out   std_logic;
          sample_out_rot_s_3   : out   std_logic;
          sample_out_rot_s_4   : out   std_logic;
          HRESETn_c            : in    std_logic;
          HCLK_c               : in    std_logic
        );

end IIR_CEL_CTRLR_v2_CONTROL;

architecture DEF_ARCH of IIR_CEL_CTRLR_v2_CONTROL is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \Chanel_ongoing_RNISG5D[13]_net_1\, 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_7, N_270, 
        Chanel_ongoing_n20, \Chanel_ongoing[20]_net_1\, N_278, 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Chanel_ongoing_n21, 
        \Chanel_ongoing[21]_net_1\, N_279, Chanel_ongoing_n22, 
        \Chanel_ongoing[22]_net_1\, N_725, Chanel_ongoing_n28, 
        \Chanel_ongoing[28]_net_1\, N_293, 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Chanel_ongoing_n29, 
        \Chanel_ongoing[29]_net_1\, N_295, Chanel_ongoing_n30, 
        \Chanel_ongoing[30]_net_1\, N_327, Chanel_ongoing_n31, 
        \Chanel_ongoing[31]_net_1\, N_335, N_250, 
        \Chanel_ongoing[0]_net_1\, \Chanel_ongoing[1]_net_1\, 
        \Chanel_ongoing[2]_net_1\, N_256, 
        \Chanel_ongoing[7]_net_1\, N_254, 
        \Chanel_ongoing[8]_net_1\, N_265, 
        \Chanel_ongoing[11]_net_1\, N_258, 
        \Chanel_ongoing[12]_net_1\, \Chanel_ongoing[13]_net_1\, 
        N_271, \Chanel_ongoing[14]_net_1\, N_272, 
        \Chanel_ongoing[15]_net_1\, N_273, 
        \Chanel_ongoing[16]_net_1\, N_275, 
        \Chanel_ongoing[17]_net_1\, N_276, 
        \Chanel_ongoing[18]_net_1\, \Chanel_ongoing[19]_net_1\, 
        N_288, \Chanel_ongoing[23]_net_1\, N_290, 
        \Chanel_ongoing[24]_net_1\, N_292, N_291, 
        \Chanel_ongoing[26]_net_1\, \Chanel_ongoing[27]_net_1\, 
        \Chanel_ongoing[9]_net_1\, \Chanel_ongoing[10]_net_1\, 
        \Chanel_ongoing[25]_net_1\, \Chanel_ongoing[5]_net_1\, 
        N_252, \Chanel_ongoing[6]_net_1\, 
        \Chanel_ongoing[3]_net_1\, \Chanel_ongoing[4]_net_1\, 
        N_75, \Cel_ongoing[29]_net_1\, \Cel_ongoing[30]_net_1\, 
        N_72, I129_un1_Y, \Cel_ongoing[13]_net_1\, N_28_0, 
        ADD_32x32_fast_I129_un1_Y_14, N_20_0, 
        \Cel_ongoing[3]_net_1\, N_18_0, \Cel_ongoing[4]_net_1\, 
        N_22_0, \Cel_ongoing[5]_net_1\, \Cel_ongoing[6]_net_1\, 
        N_24_0, \Cel_ongoing[7]_net_1\, \Cel_ongoing[8]_net_1\, 
        N_26_0, \Cel_ongoing[9]_net_1\, \Cel_ongoing[10]_net_1\, 
        \Cel_ongoing[11]_net_1\, \Cel_ongoing[12]_net_1\, N_44, 
        \Cel_ongoing[14]_net_1\, N_47, \Cel_ongoing[15]_net_1\, 
        \Cel_ongoing[16]_net_1\, N_48, N_51, 
        \Cel_ongoing[17]_net_1\, \Cel_ongoing[18]_net_1\, N_52, 
        N_55, \Cel_ongoing[19]_net_1\, \Cel_ongoing[20]_net_1\, 
        N_56, N_59, \Cel_ongoing[21]_net_1\, 
        \Cel_ongoing[22]_net_1\, N_60, N_63, 
        \Cel_ongoing[23]_net_1\, \Cel_ongoing[24]_net_1\, N_64, 
        N_66, \Cel_ongoing[25]_net_1\, N_68, 
        \Cel_ongoing[26]_net_1\, N_70, \Cel_ongoing[27]_net_1\, 
        \Cel_ongoing[28]_net_1\, \un1_IIR_CEL_STATE_17_i[17]\, 
        \Cel_ongoing_RNO[14]_net_1\, N_371_0, 
        \Cel_ongoing_RNO[15]_net_1\, N_435, N_436, N_437, N_438, 
        N_439, N_440, N_371, N_441, N_442, N_443, N_444, N_445, 
        N_446, N_447, N_448, N_449, N_450, 
        \Cel_ongoing[31]_net_1\, \Cel_ongoing[1]_net_1\, N_16_0, 
        \Cel_ongoing[2]_net_1\, \Cel_ongoing[0]_net_1\, N_566, 
        N_6, \IIR_CEL_STATE[4]_net_1\, \IIR_CEL_STATE_i[9]_net_1\, 
        \IIR_CEL_STATE[0]_net_1\, \IIR_CEL_STATE[1]_net_1\, 
        alu_selected_coeff_n0, alu_selected_coeffe, N_713, 
        N_567_i_0, \IIR_CEL_STATE[8]_net_1\, N_127_0, N_274, 
        un1_alu_sel_input_0_sqmuxa_2_i_0_s_0_0, N_452, N_248, 
        \sample_in_rot_RNI6EV7\, \IIR_CEL_STATE_i_i[9]\, 
        ADD_32x32_fast_I129_un1_Y_9, ADD_32x32_fast_I129_un1_Y_8, 
        ADD_32x32_fast_I129_un1_Y_13, ADD_32x32_fast_I129_un1_Y_5, 
        ADD_32x32_fast_I129_un1_Y_4, ADD_32x32_fast_I129_un1_Y_11, 
        ADD_32x32_fast_I129_un1_Y_7, ADD_32x32_fast_I129_un1_Y_3, 
        ADD_32x32_fast_I129_un1_Y_1, 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_2, 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_1, 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_6, 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_4, 
        Chanel_ongoing_n2_0_i_0_0, Chanel_ongoing_n7_0_i_0_0, 
        Chanel_ongoing_n6_0_i_0_0, Chanel_ongoing_n4_0_i_0_0, 
        Chanel_ongoing_n8_0_i_0_0, Chanel_ongoing_n5_0_i_0_0, 
        Chanel_ongoing_n1_0_i_0_0, alu_selected_coeff_n3_0_i_0, 
        N_717, N_733_1, N_294, N_453, alu_selected_coeff_n2_0_i_0, 
        \alu_sel_coeff_0[2]\, \Cel_ongoing_6_i_i_1[0]\, 
        \Cel_ongoing_6_i_i_a2_0_0[0]\, N_328, 
        \Cel_ongoing_6_i_i_0[0]\, 
        \un1_IIR_CEL_STATE_17_i_1_i_0[31]\, N_457, 
        un1_IIR_CEL_STATE_22_0_0, \IIR_CEL_STATE[5]_net_1\, 
        raddr_add1_2_i_a2_0_0, \IIR_CEL_STATE[3]_net_1\, 
        \in_sel_src_8_i_a2_0_a2_0_0[1]\, \IIR_CEL_STATE[6]_net_1\, 
        \IIR_CEL_STATE[7]_net_1\, Cel_ongoing_0_sqmuxa_0_a2_0_27, 
        Cel_ongoing_0_sqmuxa_0_a2_0_16, 
        Cel_ongoing_0_sqmuxa_0_a2_0_15, 
        Cel_ongoing_0_sqmuxa_0_a2_0_24, 
        Cel_ongoing_0_sqmuxa_0_a2_0_26, 
        Cel_ongoing_0_sqmuxa_0_a2_0_12, 
        Cel_ongoing_0_sqmuxa_0_a2_0_11, 
        Cel_ongoing_0_sqmuxa_0_a2_0_22, 
        Cel_ongoing_0_sqmuxa_0_a2_0_25, 
        Cel_ongoing_0_sqmuxa_0_a2_0_8, 
        Cel_ongoing_0_sqmuxa_0_a2_0_7, 
        Cel_ongoing_0_sqmuxa_0_a2_0_20, N_479, 
        Cel_ongoing_0_sqmuxa_0_a2_0_4, 
        Cel_ongoing_0_sqmuxa_0_a2_0_18, 
        Cel_ongoing_0_sqmuxa_0_a2_0_14, 
        Cel_ongoing_0_sqmuxa_0_a2_0_10, 
        Cel_ongoing_0_sqmuxa_0_a2_0_6, 
        Cel_ongoing_0_sqmuxa_0_a2_0_3, 
        Cel_ongoing_0_sqmuxa_0_a2_0_1, 
        \in_sel_src_8_i_a2_0_o2_0_27[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_18[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_17[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_23[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_26[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_12[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_11[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_22[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_25[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_8[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_7[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_20[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_2[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_1[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_15[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_14[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_10[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_6[1]\, 
        \in_sel_src_8_i_a2_0_o2_0_4[1]\, ram_write_2_0_a2_0, N_18, 
        N_20, N_650, N_651, N_703, N_206, N_480, 
        un1_IIR_CEL_STATE_20, N_325_i, N_714, 
        un1_IIR_CEL_STATE_22, N_796_i, N_736, N_723_i_0, N_737, 
        N_735, N_289, N_11, N_22, N_216, N_216_tz, N_33_0, N_34_0, 
        N_35_0, N_36_0, N_38, N_40, N_42, Chanel_ongoing_n0, 
        \Cel_ongoing_RNO[3]_net_1\, \Cel_ongoing_RNO[4]_net_1\, 
        \Cel_ongoing_RNO[5]_net_1\, \Cel_ongoing_RNO[6]_net_1\, 
        \Cel_ongoing_RNO[7]_net_1\, \Cel_ongoing_RNO[8]_net_1\, 
        \Cel_ongoing_RNO[9]_net_1\, \Cel_ongoing_RNO[10]_net_1\, 
        \Cel_ongoing_RNO[11]_net_1\, \Cel_ongoing_RNO[12]_net_1\, 
        N_462, N_374_i, N_269, N_332, Chanel_ongoing_n17, 
        Chanel_ongoing_n18, Chanel_ongoing_n19, 
        Chanel_ongoing_n23, Chanel_ongoing_n24, 
        Chanel_ongoing_n26, Chanel_ongoing_n27, N_224, N_724, 
        N_229, N_232, sample_in_rotate, N_373_i, N_372_i, N_127, 
        N_461, N_460, \IIR_CEL_STATE_ns[8]\, N_336_i_i_0, N_221, 
        \Cel_ongoing_RNO[13]_net_1\, \Cel_ongoing_RNO[1]_net_1\, 
        N_31_0, N_32_0_i_0, N_715, N_15_i, \alu_sel_coeff[3]\, 
        N_353, N_712, \IIR_CEL_STATE[2]_net_1\, N_227, N_729, 
        N_523, N_568_i_0, ram_write_2, un1_IIR_CEL_STATE_27, 
        N_477, N_569, N_334, N_180, N_204, Chanel_ongoing_n25, 
        un1_IIR_CEL_STATE_25, N_268_i_0, alu_sel_input_1, 
        sample_in_rot_2, N_512_i_0, \alu_sel_coeff[0]\, 
        \alu_sel_coeff[2]\, \alu_sel_coeff[4]\, ram_write_net_1, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    alu_sel_coeff(4) <= \alu_sel_coeff[4]\;
    alu_sel_coeff(3) <= \alu_sel_coeff[3]\;
    alu_sel_coeff(2) <= \alu_sel_coeff[2]\;
    alu_sel_coeff(0) <= \alu_sel_coeff[0]\;
    alu_sel_coeff_0_2 <= \alu_sel_coeff_0[2]\;
    ram_write <= ram_write_net_1;

    sample_in_rot_RNO : NOR2A
      port map(A => \IIR_CEL_STATE[7]_net_1\, B => N_328, Y => 
        sample_in_rot_2);
    
    \Cel_ongoing_RNIP2TO[8]\ : NOR3A
      port map(A => \in_sel_src_8_i_a2_0_o2_0_4[1]\, B => 
        \Cel_ongoing[8]_net_1\, C => \Cel_ongoing[7]_net_1\, Y
         => \in_sel_src_8_i_a2_0_o2_0_17[1]\);
    
    un1_IIR_CEL_STATE_17_m17 : NOR3C
      port map(A => \Cel_ongoing[1]_net_1\, B => N_16_0, C => 
        \Cel_ongoing[2]_net_1\, Y => N_18_0);
    
    \IIR_CEL_STATE_RNIU1T5[5]\ : OR2
      port map(A => \IIR_CEL_STATE[7]_net_1\, B => 
        \IIR_CEL_STATE[5]_net_1\, Y => N_289);
    
    \Cel_ongoing_RNO[9]\ : XA1
      port map(A => \Cel_ongoing[9]_net_1\, B => N_24_0, C => 
        N_371_0, Y => \Cel_ongoing_RNO[9]_net_1\);
    
    \in_sel_src[0]\ : DFN1E0C0
      port map(D => N_268_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => un1_IIR_CEL_STATE_27, Q => in_sel_src(0));
    
    \Chanel_ongoing_RNIFMU9[17]\ : NOR2A
      port map(A => \Chanel_ongoing[17]_net_1\, B => N_273, Y => 
        N_275);
    
    \Chanel_ongoing[1]\ : DFN1E1C0
      port map(D => N_18, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[1]_net_1\);
    
    \in_sel_src_RNO_0[1]\ : OR2
      port map(A => \IIR_CEL_STATE[6]_net_1\, B => 
        \IIR_CEL_STATE[7]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_a2_0_0[1]\);
    
    \Chanel_ongoing_RNI3OA4[8]\ : NOR3C
      port map(A => \Chanel_ongoing[7]_net_1\, B => N_254, C => 
        \Chanel_ongoing[8]_net_1\, Y => N_256);
    
    \Chanel_ongoing_RNIO3D1[2]\ : OR3C
      port map(A => \Chanel_ongoing[0]_net_1\, B => 
        \Chanel_ongoing[1]_net_1\, C => \Chanel_ongoing[2]_net_1\, 
        Y => N_250);
    
    \Cel_ongoing[23]\ : DFN1C0
      port map(D => N_442, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[23]_net_1\);
    
    \Cel_ongoing[22]\ : DFN1C0
      port map(D => N_441, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[22]_net_1\);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_7 : NOR2B
      port map(A => \Cel_ongoing[28]_net_1\, B => 
        \Cel_ongoing[29]_net_1\, Y => ADD_32x32_fast_I129_un1_Y_7);
    
    \Chanel_ongoing_RNO_0[22]\ : OR2A
      port map(A => \Chanel_ongoing[21]_net_1\, B => N_279, Y => 
        N_725);
    
    \Chanel_ongoing[29]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n29, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[29]_net_1\);
    
    \Cel_ongoing_RNO[17]\ : XA1
      port map(A => \Cel_ongoing[17]_net_1\, B => N_48, C => 
        N_371_0, Y => N_436);
    
    \Chanel_ongoing_RNIPNC7[13]\ : OR2A
      port map(A => \Chanel_ongoing[13]_net_1\, B => N_265, Y => 
        N_270);
    
    \Chanel_ongoing_RNIIB91[29]\ : NOR2
      port map(A => \Chanel_ongoing[29]_net_1\, B => 
        \Chanel_ongoing[30]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_10);
    
    \IIR_CEL_STATE_i_RNILN7F[9]\ : AOI1B
      port map(A => N_733_1, B => N_294, C => N_453, Y => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_s_0_0);
    
    \Cel_ongoing[15]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[15]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[15]_net_1\);
    
    \Cel_ongoing_RNO[16]\ : NOR2A
      port map(A => N_371_0, B => N_47, Y => N_435);
    
    \Chanel_ongoing_RNO[30]\ : XA1C
      port map(A => \Chanel_ongoing[30]_net_1\, B => N_327, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n30);
    
    \Cel_ongoing_RNO[21]\ : XA1
      port map(A => \Cel_ongoing[21]_net_1\, B => N_56, C => 
        N_371, Y => N_440);
    
    \alu_selected_coeff[4]\ : DFN1E1C0
      port map(D => N_715, CLK => HCLK_c, CLR => HRESETn_c, E => 
        alu_selected_coeffe, Q => \alu_sel_coeff[4]\);
    
    \Cel_ongoing[2]\ : DFN1C0
      port map(D => N_227, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[2]_net_1\);
    
    \alu_selected_coeff_RNIH4TI5[0]\ : NOR2A
      port map(A => N_371, B => \alu_sel_coeff[0]\, Y => 
        alu_selected_coeff_n0);
    
    \Cel_ongoing_RNIT33B[0]\ : NOR2A
      port map(A => \Cel_ongoing[0]_net_1\, B => 
        \Cel_ongoing[14]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_7[1]\);
    
    \alu_selected_coeff_RNO[3]\ : NOR2A
      port map(A => N_371_0, B => alu_selected_coeff_n3_0_i_0, Y
         => N_714);
    
    \Chanel_ongoing_RNO_0[9]\ : XNOR2
      port map(A => N_256, B => \Chanel_ongoing[9]_net_1\, Y => 
        N_372_i);
    
    \IIR_CEL_STATE_RNO[2]\ : NOR2A
      port map(A => \IIR_CEL_STATE[4]_net_1\, B => N_523, Y => 
        N_477);
    
    \Chanel_ongoing_RNIQVNF[26]\ : OR2B
      port map(A => N_291, B => \Chanel_ongoing[26]_net_1\, Y => 
        N_292);
    
    alu_sel_input_RNO : NOR2
      port map(A => \IIR_CEL_STATE[6]_net_1\, B => 
        \IIR_CEL_STATE[4]_net_1\, Y => alu_sel_input_1);
    
    \Chanel_ongoing_RNO_0[3]\ : XNOR2
      port map(A => N_250, B => \Chanel_ongoing[3]_net_1\, Y => 
        N_336_i_i_0);
    
    \Cel_ongoing_RNO_1[0]\ : NOR2B
      port map(A => \IIR_CEL_STATE[4]_net_1\, B => 
        \un1_IIR_CEL_STATE_17_i_1_i_0[31]\, Y => 
        \Cel_ongoing_6_i_i_a2_0_0[0]\);
    
    \Chanel_ongoing[30]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n30, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[30]_net_1\);
    
    \IIR_CEL_STATE_RNI5V1J5[2]\ : OR2B
      port map(A => N_371, B => N_353, Y => alu_selected_coeffe);
    
    \Cel_ongoing_RNO[5]\ : NOR2A
      port map(A => N_371_0, B => N_35_0, Y => 
        \Cel_ongoing_RNO[5]_net_1\);
    
    \Cel_ongoing_RNIDJOG[18]\ : NOR3A
      port map(A => \in_sel_src_8_i_a2_0_o2_0_10[1]\, B => 
        \Cel_ongoing[18]_net_1\, C => \Cel_ongoing[17]_net_1\, Y
         => \in_sel_src_8_i_a2_0_o2_0_20[1]\);
    
    \Cel_ongoing[24]\ : DFN1C0
      port map(D => N_443, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[24]_net_1\);
    
    un1_IIR_CEL_STATE_17_m54 : AX1E
      port map(A => \Cel_ongoing[19]_net_1\, B => N_52, C => 
        \Cel_ongoing[20]_net_1\, Y => N_55);
    
    \Chanel_ongoing_RNIDQB2[4]\ : NOR3B
      port map(A => \Chanel_ongoing[3]_net_1\, B => 
        \Chanel_ongoing[4]_net_1\, C => N_250, Y => N_252);
    
    \IIR_CEL_STATE_i[9]\ : DFN1
      port map(D => N_512_i_0, CLK => HCLK_c, Q => 
        \IIR_CEL_STATE_i[9]_net_1\);
    
    \Chanel_ongoing_RNI61B3[6]\ : NOR3C
      port map(A => \Chanel_ongoing[5]_net_1\, B => N_252, C => 
        \Chanel_ongoing[6]_net_1\, Y => N_254);
    
    \Chanel_ongoing[8]\ : DFN1E1C0
      port map(D => N_651, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[8]_net_1\);
    
    \Chanel_ongoing_RNO[13]\ : XA1C
      port map(A => \Chanel_ongoing[13]_net_1\, B => N_265, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => N_224);
    
    \Chanel_ongoing_RNIKIU[2]\ : NOR2
      port map(A => \Chanel_ongoing[2]_net_1\, B => 
        \Chanel_ongoing[4]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_1);
    
    \Cel_ongoing_RNO[11]\ : XA1
      port map(A => \Cel_ongoing[11]_net_1\, B => N_26_0, C => 
        N_371_0, Y => \Cel_ongoing_RNO[11]_net_1\);
    
    \Cel_ongoing_RNIKMF11[22]\ : NOR3C
      port map(A => \in_sel_src_8_i_a2_0_o2_0_12[1]\, B => 
        \in_sel_src_8_i_a2_0_o2_0_11[1]\, C => 
        \in_sel_src_8_i_a2_0_o2_0_22[1]\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_26[1]\);
    
    \IIR_CEL_STATE_RNIRIR8[6]\ : OR3
      port map(A => \IIR_CEL_STATE[3]_net_1\, B => 
        \IIR_CEL_STATE[6]_net_1\, C => \IIR_CEL_STATE[7]_net_1\, 
        Y => N_334);
    
    \alu_selected_coeff_RNO_0[4]\ : AX1A
      port map(A => N_717, B => \alu_sel_coeff[3]\, C => 
        \alu_sel_coeff[4]\, Y => N_15_i);
    
    \Chanel_ongoing[3]\ : DFN1E1C0
      port map(D => N_221, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[3]_net_1\);
    
    \Chanel_ongoing_RNO_0[6]\ : AX1E
      port map(A => \Chanel_ongoing[5]_net_1\, B => N_252, C => 
        \Chanel_ongoing[6]_net_1\, Y => Chanel_ongoing_n6_0_i_0_0);
    
    ram_write_RNO : AO1B
      port map(A => ram_write_2_0_a2_0, B => N_733_1, C => N_480, 
        Y => ram_write_2);
    
    \Cel_ongoing_RNICE615_0[2]\ : OR2A
      port map(A => N_325_i, B => \Cel_ongoing[2]_net_1\, Y => 
        N_332);
    
    \Cel_ongoing[0]\ : DFN1C0
      port map(D => N_206, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[0]_net_1\);
    
    sample_out_rot_3 : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s_3);
    
    \IIR_CEL_STATE_RNISQ2Q5[2]\ : AO1
      port map(A => N_523, B => \IIR_CEL_STATE[4]_net_1\, C => 
        \IIR_CEL_STATE[2]_net_1\, Y => un1_IIR_CEL_STATE_27);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_13 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_5, B => 
        ADD_32x32_fast_I129_un1_Y_4, C => 
        ADD_32x32_fast_I129_un1_Y_11, Y => 
        ADD_32x32_fast_I129_un1_Y_13);
    
    \Chanel_ongoing_RNIE545[14]\ : NOR3C
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_12, B => 
        Cel_ongoing_0_sqmuxa_0_a2_0_11, C => 
        Cel_ongoing_0_sqmuxa_0_a2_0_22, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_26);
    
    \IIR_CEL_STATE_RNI9V445[4]\ : OR2B
      port map(A => N_328, B => \IIR_CEL_STATE[4]_net_1\, Y => 
        N_248);
    
    \IIR_CEL_STATE_i_RNILP76[9]\ : OR3
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => 
        sample_val_delay, C => \IIR_CEL_STATE[4]_net_1\, Y => 
        N_453);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_4 : NOR2B
      port map(A => \Cel_ongoing[22]_net_1\, B => 
        \Cel_ongoing[23]_net_1\, Y => ADD_32x32_fast_I129_un1_Y_4);
    
    un1_IIR_CEL_STATE_17_m50 : AX1E
      port map(A => \Cel_ongoing[17]_net_1\, B => N_48, C => 
        \Cel_ongoing[18]_net_1\, Y => N_51);
    
    \IIR_CEL_STATE_i_RNIEAL96[9]\ : OR2B
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0_s_0_0, B => 
        N_452, Y => un1_alu_sel_input_0_sqmuxa_2_i_0_0);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y : NOR3C
      port map(A => \Cel_ongoing[13]_net_1\, B => N_28_0, C => 
        ADD_32x32_fast_I129_un1_Y_14, Y => I129_un1_Y);
    
    \IIR_CEL_STATE[2]\ : DFN1E1
      port map(D => N_477, CLK => HCLK_c, E => HRESETn_c, Q => 
        \IIR_CEL_STATE[2]_net_1\);
    
    \Chanel_ongoing[13]\ : DFN1E1C0
      port map(D => N_224, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[13]_net_1\);
    
    \Chanel_ongoing[12]\ : DFN1E1C0
      port map(D => N_216, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[12]_net_1\);
    
    ram_write_RNO_0 : NOR2
      port map(A => \IIR_CEL_STATE[3]_net_1\, B => 
        \IIR_CEL_STATE[7]_net_1\, Y => ram_write_2_0_a2_0);
    
    un1_IIR_CEL_STATE_17_m34 : XNOR2
      port map(A => N_20_0, B => \Cel_ongoing[5]_net_1\, Y => 
        N_35_0);
    
    \IIR_CEL_STATE_i_RNIEAL96_0[9]\ : OR2B
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0_s_0_0, B => 
        N_452, Y => un1_alu_sel_input_0_sqmuxa_2_i_0);
    
    \Cel_ongoing_RNO_0[0]\ : AOI1B
      port map(A => \Cel_ongoing_6_i_i_a2_0_0[0]\, B => N_328, C
         => \Cel_ongoing_6_i_i_0[0]\, Y => 
        \Cel_ongoing_6_i_i_1[0]\);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_8 : NOR3C
      port map(A => \Cel_ongoing[15]_net_1\, B => 
        \Cel_ongoing[14]_net_1\, C => ADD_32x32_fast_I129_un1_Y_1, 
        Y => ADD_32x32_fast_I129_un1_Y_8);
    
    sample_out_rot_1 : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s_1);
    
    \Chanel_ongoing_RNI9OEE[24]\ : OR2A
      port map(A => \Chanel_ongoing[24]_net_1\, B => N_288, Y => 
        N_290);
    
    \Cel_ongoing_RNO[31]\ : XA1
      port map(A => \Cel_ongoing[31]_net_1\, B => N_75, C => 
        N_371, Y => N_450);
    
    \Cel_ongoing_RNIRLC8[27]\ : NOR2
      port map(A => \Cel_ongoing[27]_net_1\, B => 
        \Cel_ongoing[28]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_14[1]\);
    
    \Chanel_ongoing_RNO[31]\ : XA1C
      port map(A => \Chanel_ongoing[31]_net_1\, B => N_335, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n31);
    
    \Chanel_ongoing_RNIH791[25]\ : NOR2
      port map(A => \Chanel_ongoing[25]_net_1\, B => 
        \Chanel_ongoing[26]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_8);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_11 : NOR3C
      port map(A => \Cel_ongoing[27]_net_1\, B => 
        \Cel_ongoing[26]_net_1\, C => ADD_32x32_fast_I129_un1_Y_7, 
        Y => ADD_32x32_fast_I129_un1_Y_11);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_14 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_9, B => 
        ADD_32x32_fast_I129_un1_Y_8, C => 
        ADD_32x32_fast_I129_un1_Y_13, Y => 
        ADD_32x32_fast_I129_un1_Y_14);
    
    \Chanel_ongoing[11]\ : DFN1E1C0
      port map(D => N_462, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[11]_net_1\);
    
    \IIR_CEL_STATE[4]\ : DFN1E1
      port map(D => \IIR_CEL_STATE[3]_net_1\, CLK => HCLK_c, E
         => HRESETn_c, Q => \IIR_CEL_STATE[4]_net_1\);
    
    \Chanel_ongoing_RNI3PO5[15]\ : NOR3C
      port map(A => Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_2, B => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_1, C => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_6, Y => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_7);
    
    un1_IIR_CEL_STATE_17_m21 : NOR3C
      port map(A => \Cel_ongoing[5]_net_1\, B => N_20_0, C => 
        \Cel_ongoing[6]_net_1\, Y => N_22_0);
    
    \IIR_CEL_STATE_i_RNI16EG5[9]\ : OR2A
      port map(A => N_371, B => N_274, Y => N_127_0);
    
    \alu_selected_coeff_RNO[1]\ : NOR2B
      port map(A => S_i_0(33), B => N_371, Y => N_712);
    
    \IIR_CEL_STATE_RNI3D16[1]\ : NOR3A
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => 
        \IIR_CEL_STATE[0]_net_1\, C => \IIR_CEL_STATE[1]_net_1\, 
        Y => N_6);
    
    \Cel_ongoing_RNIJEQD[6]\ : NOR2
      port map(A => \Cel_ongoing[5]_net_1\, B => 
        \Cel_ongoing[6]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_2[1]\);
    
    un1_IIR_CEL_STATE_17_m30 : XNOR2
      port map(A => N_16_0, B => \Cel_ongoing[1]_net_1\, Y => 
        N_31_0);
    
    \Chanel_ongoing_RNO[20]\ : XA1C
      port map(A => \Chanel_ongoing[20]_net_1\, B => N_278, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n20);
    
    \Chanel_ongoing[20]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n20, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[20]_net_1\);
    
    \Chanel_ongoing_RNIUQV[7]\ : NOR2
      port map(A => \Chanel_ongoing[7]_net_1\, B => 
        \Chanel_ongoing[9]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_3);
    
    \Chanel_ongoing_RNIFUT[1]\ : NOR2
      port map(A => \Chanel_ongoing[1]_net_1\, B => 
        \Chanel_ongoing[0]_net_1\, Y => N_479);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Chanel_ongoing[27]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n27, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[27]_net_1\);
    
    \Cel_ongoing_RNO[25]\ : XA1
      port map(A => \Cel_ongoing[25]_net_1\, B => N_64, C => 
        N_371, Y => N_444);
    
    \Chanel_ongoing_RNO_0[7]\ : XOR2
      port map(A => \Chanel_ongoing[7]_net_1\, B => N_254, Y => 
        Chanel_ongoing_n7_0_i_0_0);
    
    un1_IIR_CEL_STATE_17_m71 : NOR2B
      port map(A => N_70, B => \Cel_ongoing[28]_net_1\, Y => N_72);
    
    \Chanel_ongoing_RNII4QD[23]\ : OR2A
      port map(A => \Chanel_ongoing[23]_net_1\, B => 
        \Chanel_ongoing_RNISG5D[13]_net_1\, Y => N_288);
    
    \alu_selected_coeff_RNIR19H[2]\ : OR2A
      port map(A => \alu_sel_coeff[2]\, B => S(8), Y => N_717);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    raddr_add1_RNO_0 : OR3
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => 
        sample_val_delay, C => \IIR_CEL_STATE[3]_net_1\, Y => 
        N_737);
    
    \Chanel_ongoing_RNO_0[12]\ : AX1E
      port map(A => \Chanel_ongoing[11]_net_1\, B => N_258, C => 
        \Chanel_ongoing[12]_net_1\, Y => N_216_tz);
    
    \Chanel_ongoing_RNI9Q63[19]\ : NOR3C
      port map(A => \Chanel_ongoing[20]_net_1\, B => 
        \Chanel_ongoing[19]_net_1\, C => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_4, Y => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_6);
    
    sample_out_rot_0 : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s_0);
    
    \Chanel_ongoing_RNIF71H[28]\ : OR2A
      port map(A => \Chanel_ongoing[28]_net_1\, B => N_293, Y => 
        N_295);
    
    \IIR_CEL_STATE[5]\ : DFN1E1
      port map(D => N_204, CLK => HCLK_c, E => HRESETn_c, Q => 
        \IIR_CEL_STATE[5]_net_1\);
    
    \Cel_ongoing[25]\ : DFN1C0
      port map(D => N_444, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[25]_net_1\);
    
    \IIR_CEL_STATE_RNO[5]\ : OR2A
      port map(A => N_248, B => N_353, Y => N_204);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_5 : NOR2B
      port map(A => \Cel_ongoing[24]_net_1\, B => 
        \Cel_ongoing[25]_net_1\, Y => ADD_32x32_fast_I129_un1_Y_5);
    
    \Chanel_ongoing[18]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n18, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[18]_net_1\);
    
    \Chanel_ongoing[16]\ : DFN1E1C0
      port map(D => N_232, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[16]_net_1\);
    
    \alu_selected_coeff[3]\ : DFN1E1C0
      port map(D => N_714, CLK => HCLK_c, CLR => HRESETn_c, E => 
        alu_selected_coeffe, Q => \alu_sel_coeff[3]\);
    
    \Chanel_ongoing_RNITMT1[22]\ : NOR3C
      port map(A => \Chanel_ongoing[14]_net_1\, B => 
        \Chanel_ongoing[22]_net_1\, C => 
        \Chanel_ongoing[21]_net_1\, Y => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_4);
    
    \Cel_ongoing_RNO[15]\ : XA1
      port map(A => \Cel_ongoing[15]_net_1\, B => N_44, C => 
        N_371_0, Y => \Cel_ongoing_RNO[15]_net_1\);
    
    un1_IIR_CEL_STATE_17_m67 : NOR2B
      port map(A => N_66, B => \Cel_ongoing[26]_net_1\, Y => N_68);
    
    \alu_ctrl[0]\ : DFN1E0C0
      port map(D => N_568_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[2]_net_1\, Q => alu_ctrl(0));
    
    raddr_add1_RNO_1 : OR3B
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => N_289, C => 
        \IIR_CEL_STATE[3]_net_1\, Y => N_735);
    
    \Chanel_ongoing_RNI7791[20]\ : NOR2
      port map(A => \Chanel_ongoing[20]_net_1\, B => 
        \Chanel_ongoing[21]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_14);
    
    \Cel_ongoing_RNIU5UA1[31]\ : NOR3C
      port map(A => \in_sel_src_8_i_a2_0_o2_0_2[1]\, B => 
        \in_sel_src_8_i_a2_0_o2_0_1[1]\, C => 
        \in_sel_src_8_i_a2_0_o2_0_15[1]\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_23[1]\);
    
    un1_IIR_CEL_STATE_17_m23 : NOR3C
      port map(A => \Cel_ongoing[7]_net_1\, B => N_22_0, C => 
        \Cel_ongoing[8]_net_1\, Y => N_24_0);
    
    \Chanel_ongoing_RNI2NL8[15]\ : OR2A
      port map(A => \Chanel_ongoing[15]_net_1\, B => N_271, Y => 
        N_272);
    
    \Chanel_ongoing[14]\ : DFN1E1C0
      port map(D => N_724, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[14]_net_1\);
    
    \IIR_CEL_STATE_i_RNIO893[9]\ : NOR2A
      port map(A => sample_val_delay, B => 
        \IIR_CEL_STATE_i[9]_net_1\, Y => N_274);
    
    \alu_ctrl[2]\ : DFN1E0C0
      port map(D => \IIR_CEL_STATE_i_i[9]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \IIR_CEL_STATE[2]_net_1\, Q => 
        alu_ctrl(2));
    
    \Chanel_ongoing_RNO[10]\ : NOR2
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0, B => 
        N_373_i, Y => N_461);
    
    \ram_sel_Wdata[1]\ : DFN1E0C0
      port map(D => un1_IIR_CEL_STATE_22, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \IIR_CEL_STATE[8]_net_1\, Q => 
        ram_sel_Wdata(1));
    
    \IIR_CEL_STATE_RNIN1T5[5]\ : NOR2
      port map(A => \IIR_CEL_STATE[0]_net_1\, B => 
        \IIR_CEL_STATE[5]_net_1\, Y => un1_IIR_CEL_STATE_22_0_0);
    
    \Chanel_ongoing_RNIBV81[15]\ : NOR2B
      port map(A => \Chanel_ongoing[15]_net_1\, B => 
        \Chanel_ongoing[16]_net_1\, Y => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_1);
    
    \Cel_ongoing_RNO[4]\ : NOR2A
      port map(A => N_371_0, B => N_34_0, Y => 
        \Cel_ongoing_RNO[4]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Chanel_ongoing_RNO_0[11]\ : XNOR2
      port map(A => N_258, B => \Chanel_ongoing[11]_net_1\, Y => 
        N_374_i);
    
    \Chanel_ongoing_RNID791[23]\ : NOR2
      port map(A => \Chanel_ongoing[23]_net_1\, B => 
        \Chanel_ongoing[24]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_7);
    
    \Cel_ongoing[4]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[4]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[4]_net_1\);
    
    \Chanel_ongoing_RNO[21]\ : XA1C
      port map(A => \Chanel_ongoing[21]_net_1\, B => N_279, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n21);
    
    \Chanel_ongoing_RNI76JA[18]\ : OR2B
      port map(A => N_275, B => \Chanel_ongoing[18]_net_1\, Y => 
        N_276);
    
    \Chanel_ongoing_RNO[29]\ : XA1C
      port map(A => \Chanel_ongoing[29]_net_1\, B => N_295, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n29);
    
    \Chanel_ongoing_RNIJ9SB[20]\ : OR2A
      port map(A => \Chanel_ongoing[20]_net_1\, B => N_278, Y => 
        N_279);
    
    \alu_ctrl[1]\ : DFN1E0C0
      port map(D => N_569, CLK => HCLK_c, CLR => HRESETn_c, E => 
        \IIR_CEL_STATE[2]_net_1\, Q => alu_ctrl(1));
    
    sample_out_val : DFN1E0C0
      port map(D => \IIR_CEL_STATE[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => N_353, Q => sample_out_val_s);
    
    raddr_add1_RNO_3 : OR2A
      port map(A => \IIR_CEL_STATE[3]_net_1\, B => N_274, Y => 
        raddr_add1_2_i_a2_0_0);
    
    \Chanel_ongoing[31]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n31, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[31]_net_1\);
    
    un1_IIR_CEL_STATE_17_m29 : XNOR2
      port map(A => N_566, B => \Cel_ongoing[0]_net_1\, Y => 
        \un1_IIR_CEL_STATE_17_i_1_i_0[31]\);
    
    \IIR_CEL_STATE_RNI0UV8[4]\ : NOR2A
      port map(A => N_6, B => \IIR_CEL_STATE[4]_net_1\, Y => 
        N_566);
    
    \Cel_ongoing_RNI679Q4[12]\ : NOR3C
      port map(A => \in_sel_src_8_i_a2_0_o2_0_26[1]\, B => 
        \in_sel_src_8_i_a2_0_o2_0_25[1]\, C => 
        \in_sel_src_8_i_a2_0_o2_0_27[1]\, Y => N_325_i);
    
    sample_out_rot_2 : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s_2);
    
    \Chanel_ongoing_RNI53M8[6]\ : NOR3C
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_16, B => 
        Cel_ongoing_0_sqmuxa_0_a2_0_15, C => 
        Cel_ongoing_0_sqmuxa_0_a2_0_24, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_27);
    
    \Chanel_ongoing_RNIO6I2[18]\ : NOR3A
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_14, B => 
        \Chanel_ongoing[19]_net_1\, C => 
        \Chanel_ongoing[18]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_22);
    
    \Chanel_ongoing_RNI1C3F[25]\ : NOR2A
      port map(A => \Chanel_ongoing[25]_net_1\, B => N_290, Y => 
        N_291);
    
    un1_IIR_CEL_STATE_17_m19 : NOR3C
      port map(A => \Cel_ongoing[3]_net_1\, B => N_18_0, C => 
        \Cel_ongoing[4]_net_1\, Y => N_20_0);
    
    \IIR_CEL_STATE_RNI9T4D5[4]\ : OR2A
      port map(A => N_248, B => N_566, Y => N_371_0);
    
    un1_IIR_CEL_STATE_17_m46 : AX1E
      port map(A => \Cel_ongoing[15]_net_1\, B => N_44, C => 
        \Cel_ongoing[16]_net_1\, Y => N_47);
    
    \Chanel_ongoing_RNIKJCG[27]\ : OR2A
      port map(A => \Chanel_ongoing[27]_net_1\, B => N_292, Y => 
        N_293);
    
    \Chanel_ongoing_RNI39F5[10]\ : NOR3C
      port map(A => \Chanel_ongoing[9]_net_1\, B => N_256, C => 
        \Chanel_ongoing[10]_net_1\, Y => N_258);
    
    \waddr_previous[1]\ : DFN1E0C0
      port map(D => N_729, CLK => HCLK_c, CLR => HRESETn_c, E => 
        \IIR_CEL_STATE[8]_net_1\, Q => waddr_previous(1));
    
    un1_IIR_CEL_STATE_17_m37 : AX1E
      port map(A => \Cel_ongoing[7]_net_1\, B => N_22_0, C => 
        \Cel_ongoing[8]_net_1\, Y => N_38);
    
    un1_IIR_CEL_STATE_17_m25 : NOR3C
      port map(A => \Cel_ongoing[9]_net_1\, B => N_24_0, C => 
        \Cel_ongoing[10]_net_1\, Y => N_26_0);
    
    \Cel_ongoing_RNIF5B8[22]\ : NOR2
      port map(A => \Cel_ongoing[21]_net_1\, B => 
        \Cel_ongoing[22]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_11[1]\);
    
    raddr_add1_RNO : NOR3C
      port map(A => N_737, B => N_735, C => N_736, Y => N_723_i_0);
    
    un1_IIR_CEL_STATE_17_m15 : NOR2A
      port map(A => \Cel_ongoing[0]_net_1\, B => N_566, Y => 
        N_16_0);
    
    \IIR_CEL_STATE_RNI1A4N5[4]\ : NOR2
      port map(A => N_796_i, B => N_480, Y => 
        \IIR_CEL_STATE_ns[8]\);
    
    \IIR_CEL_STATE[7]\ : DFN1E1
      port map(D => \IIR_CEL_STATE[6]_net_1\, CLK => HCLK_c, E
         => HRESETn_c, Q => \IIR_CEL_STATE[7]_net_1\);
    
    \IIR_CEL_STATE_RNIL1T5[1]\ : OR2
      port map(A => \IIR_CEL_STATE[2]_net_1\, B => 
        \IIR_CEL_STATE[1]_net_1\, Y => N_567_i_0);
    
    \Cel_ongoing[19]\ : DFN1C0
      port map(D => N_438, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[19]_net_1\);
    
    \Chanel_ongoing_RNO[11]\ : NOR2
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0_0, B => 
        N_374_i, Y => N_462);
    
    \Chanel_ongoing_RNO[24]\ : XA1C
      port map(A => \Chanel_ongoing[24]_net_1\, B => N_288, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n24);
    
    \Chanel_ongoing_RNO[19]\ : XA1C
      port map(A => \Chanel_ongoing[19]_net_1\, B => N_276, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n19);
    
    \Chanel_ongoing_RNIN1V1[6]\ : NOR3A
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_3, B => 
        \Chanel_ongoing[6]_net_1\, C => \Chanel_ongoing[5]_net_1\, 
        Y => Cel_ongoing_0_sqmuxa_0_a2_0_16);
    
    \Chanel_ongoing[15]\ : DFN1E1C0
      port map(D => N_229, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[15]_net_1\);
    
    \Cel_ongoing[31]\ : DFN1C0
      port map(D => N_450, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[31]_net_1\);
    
    \IIR_CEL_STATE_i_RNIPIDQ5[9]\ : OR2A
      port map(A => \IIR_CEL_STATE_ns[8]\, B => N_274, Y => N_452);
    
    \Cel_ongoing_RNIJLB8[24]\ : NOR2
      port map(A => \Cel_ongoing[23]_net_1\, B => 
        \Cel_ongoing[24]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_12[1]\);
    
    \alu_selected_coeff_RNO[4]\ : NOR2A
      port map(A => N_371, B => N_15_i, Y => N_715);
    
    \Cel_ongoing[30]\ : DFN1C0
      port map(D => N_449, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[30]_net_1\);
    
    \Chanel_ongoing_RNO_0[5]\ : XNOR2
      port map(A => \Chanel_ongoing[5]_net_1\, B => N_252, Y => 
        Chanel_ongoing_n5_0_i_0_0);
    
    \Chanel_ongoing[6]\ : DFN1E1C0
      port map(D => N_22, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[6]_net_1\);
    
    \alu_selected_coeff_RNO_0[3]\ : XOR2
      port map(A => N_717, B => \alu_sel_coeff[3]\, Y => 
        alu_selected_coeff_n3_0_i_0);
    
    sample_out_rot : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s);
    
    \Chanel_ongoing[23]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n23, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[23]_net_1\);
    
    \Chanel_ongoing[22]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n22, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[22]_net_1\);
    
    sample_out_rot_4 : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => sample_out_rot_s_4);
    
    \Cel_ongoing_RNO[7]\ : XA1
      port map(A => \Cel_ongoing[7]_net_1\, B => N_22_0, C => 
        N_371_0, Y => \Cel_ongoing_RNO[7]_net_1\);
    
    ram_write_RNI0IG : INV
      port map(A => ram_write_net_1, Y => ram_write_i);
    
    \IIR_CEL_STATE_RNI012A5[5]\ : OR2B
      port map(A => un1_IIR_CEL_STATE_22_0_0, B => N_480, Y => 
        un1_IIR_CEL_STATE_22);
    
    \in_sel_src_RNO[0]\ : MX2A
      port map(A => N_334, B => N_332, S => 
        \IIR_CEL_STATE[5]_net_1\, Y => N_268_i_0);
    
    \waddr_previous[0]\ : DFN1E0C0
      port map(D => un1_IIR_CEL_STATE_25, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \IIR_CEL_STATE[8]_net_1\, Q => 
        waddr_previous(0));
    
    \Chanel_ongoing_RNI68O6[12]\ : OR3C
      port map(A => \Chanel_ongoing[11]_net_1\, B => N_258, C => 
        \Chanel_ongoing[12]_net_1\, Y => N_265);
    
    \alu_selected_coeff_0[2]\ : DFN1E1C0
      port map(D => N_713, CLK => HCLK_c, CLR => HRESETn_c, E => 
        alu_selected_coeffe, Q => \alu_sel_coeff_0[2]\);
    
    \Chanel_ongoing[21]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n21, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[21]_net_1\);
    
    \alu_selected_coeff_0[0]\ : DFN1E1C0
      port map(D => alu_selected_coeff_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => alu_selected_coeffe, Q => 
        alu_sel_coeff_0_0);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_9 : NOR3C
      port map(A => \Cel_ongoing[19]_net_1\, B => 
        \Cel_ongoing[18]_net_1\, C => ADD_32x32_fast_I129_un1_Y_3, 
        Y => ADD_32x32_fast_I129_un1_Y_9);
    
    \Cel_ongoing_RNO[22]\ : NOR2A
      port map(A => N_371, B => N_59, Y => N_441);
    
    \Chanel_ongoing_RNIDPT1[8]\ : NOR3B
      port map(A => \Chanel_ongoing[3]_net_1\, B => 
        Cel_ongoing_0_sqmuxa_0_a2_0_1, C => 
        \Chanel_ongoing[8]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_15);
    
    un1_IIR_CEL_STATE_17_m51 : NOR3C
      port map(A => \Cel_ongoing[17]_net_1\, B => N_48, C => 
        \Cel_ongoing[18]_net_1\, Y => N_52);
    
    \Chanel_ongoing_RNO[14]\ : XA1C
      port map(A => \Chanel_ongoing[14]_net_1\, B => N_270, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => N_724);
    
    \Cel_ongoing_RNISAMG[12]\ : NOR3A
      port map(A => \in_sel_src_8_i_a2_0_o2_0_6[1]\, B => 
        \Cel_ongoing[12]_net_1\, C => \Cel_ongoing[11]_net_1\, Y
         => \in_sel_src_8_i_a2_0_o2_0_18[1]\);
    
    \Cel_ongoing_RNIKTB8[20]\ : NOR2
      port map(A => \Cel_ongoing[19]_net_1\, B => 
        \Cel_ongoing[20]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_10[1]\);
    
    \raddr_rst\ : DFN1E0C0
      port map(D => un1_IIR_CEL_STATE_20, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_353, Q => raddr_rst);
    
    \Chanel_ongoing_RNIO6A9[16]\ : OR2A
      port map(A => \Chanel_ongoing[16]_net_1\, B => N_272, Y => 
        N_273);
    
    \Cel_ongoing_RNO[3]\ : NOR2A
      port map(A => N_371_0, B => N_33_0, Y => 
        \Cel_ongoing_RNO[3]_net_1\);
    
    \Chanel_ongoing_RNI18P4[1]\ : NOR3C
      port map(A => N_479, B => Cel_ongoing_0_sqmuxa_0_a2_0_4, C
         => Cel_ongoing_0_sqmuxa_0_a2_0_18, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_24);
    
    \IIR_CEL_STATE_i_RNO[9]\ : MX2B
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => N_180, S => 
        HRESETn_c, Y => N_512_i_0);
    
    \Chanel_ongoing_RNISG5D[13]\ : OR2A
      port map(A => Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_7, B => 
        N_270, Y => \Chanel_ongoing_RNISG5D[13]_net_1\);
    
    un1_IIR_CEL_STATE_17_m47 : NOR3C
      port map(A => \Cel_ongoing[15]_net_1\, B => N_44, C => 
        \Cel_ongoing[16]_net_1\, Y => N_48);
    
    \Chanel_ongoing_RNO[26]\ : XA1B
      port map(A => \Chanel_ongoing[26]_net_1\, B => N_291, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n26);
    
    \Cel_ongoing[18]\ : DFN1C0
      port map(D => N_437, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[18]_net_1\);
    
    \alu_selected_coeff_0_RNIF4EQ5[2]\ : NOR2B
      port map(A => alu_selected_coeff_n2_0_i_0, B => N_371_0, Y
         => N_713);
    
    \Chanel_ongoing_RNIHAI2[31]\ : NOR3A
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_6, B => 
        \Chanel_ongoing[12]_net_1\, C => 
        \Chanel_ongoing[31]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_18);
    
    \Cel_ongoing_RNO[12]\ : NOR2A
      port map(A => N_371_0, B => N_42, Y => 
        \Cel_ongoing_RNO[12]_net_1\);
    
    \Cel_ongoing_RNI2K2B[10]\ : NOR2
      port map(A => \Cel_ongoing[9]_net_1\, B => 
        \Cel_ongoing[10]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_4[1]\);
    
    \alu_selected_coeff[0]\ : DFN1E1C0
      port map(D => alu_selected_coeff_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => alu_selected_coeffe, Q => 
        \alu_sel_coeff[0]\);
    
    \Chanel_ongoing[19]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n19, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[19]_net_1\);
    
    \Cel_ongoing_RNI4P5K5[2]\ : OR2A
      port map(A => N_796_i, B => N_328, Y => N_523);
    
    \Cel_ongoing[16]\ : DFN1C0
      port map(D => N_435, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[16]_net_1\);
    
    un1_IIR_CEL_STATE_17_m63 : NOR3C
      port map(A => \Cel_ongoing[23]_net_1\, B => N_60, C => 
        \Cel_ongoing[24]_net_1\, Y => N_64);
    
    \Chanel_ongoing_RNO[0]\ : NOR2
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0_0, B => 
        \Chanel_ongoing[0]_net_1\, Y => Chanel_ongoing_n0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Chanel_ongoing_RNO[25]\ : XA1C
      port map(A => \Chanel_ongoing[25]_net_1\, B => N_290, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n25);
    
    \in_sel_src_RNO[1]\ : MX2
      port map(A => \in_sel_src_8_i_a2_0_a2_0_0[1]\, B => N_289, 
        S => N_332, Y => N_269);
    
    \Cel_ongoing_RNO[23]\ : XA1
      port map(A => \Cel_ongoing[23]_net_1\, B => N_60, C => 
        N_371, Y => N_442);
    
    \Chanel_ongoing[28]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n28, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[28]_net_1\);
    
    un1_IIR_CEL_STATE_17_m31 : AX1C
      port map(A => \Cel_ongoing[1]_net_1\, B => N_16_0, C => 
        \Cel_ongoing[2]_net_1\, Y => N_32_0_i_0);
    
    \Chanel_ongoing[26]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n26, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[26]_net_1\);
    
    \Chanel_ongoing_RNO[4]\ : NOR2
      port map(A => Chanel_ongoing_n4_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_11);
    
    \Cel_ongoing_RNIF5B8[30]\ : NOR2
      port map(A => \Cel_ongoing[13]_net_1\, B => 
        \Cel_ongoing[30]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_6[1]\);
    
    \Chanel_ongoing[2]\ : DFN1E1C0
      port map(D => N_703, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[2]_net_1\);
    
    \Chanel_ongoing_RNI1V81[10]\ : NOR2
      port map(A => \Chanel_ongoing[10]_net_1\, B => 
        \Chanel_ongoing[11]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_4);
    
    \Chanel_ongoing_RNO[6]\ : NOR2
      port map(A => Chanel_ongoing_n6_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_22);
    
    \IIR_CEL_STATE[6]\ : DFN1E1
      port map(D => \IIR_CEL_STATE[5]_net_1\, CLK => HCLK_c, E
         => HRESETn_c, Q => \IIR_CEL_STATE[6]_net_1\);
    
    \Cel_ongoing[17]\ : DFN1C0
      port map(D => N_436, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[17]_net_1\);
    
    \Chanel_ongoing[24]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n24, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[24]_net_1\);
    
    \Cel_ongoing_RNO[2]\ : AO1
      port map(A => N_32_0_i_0, B => N_371, C => 
        \IIR_CEL_STATE_ns[8]\, Y => N_227);
    
    \Cel_ongoing_RNIS89F[31]\ : NOR3
      port map(A => \Cel_ongoing[1]_net_1\, B => 
        \Cel_ongoing[31]_net_1\, C => \Cel_ongoing[29]_net_1\, Y
         => \in_sel_src_8_i_a2_0_o2_0_15[1]\);
    
    \Cel_ongoing[11]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[11]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[11]_net_1\);
    
    un1_IIR_CEL_STATE_17_m62 : AX1E
      port map(A => \Cel_ongoing[23]_net_1\, B => N_60, C => 
        \Cel_ongoing[24]_net_1\, Y => N_63);
    
    \Chanel_ongoing_RNO[2]\ : NOR2A
      port map(A => Chanel_ongoing_n2_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_703);
    
    \Cel_ongoing[10]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[10]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[10]_net_1\);
    
    \IIR_CEL_STATE_i_RNI16EG5_0[9]\ : OR2A
      port map(A => N_371, B => N_274, Y => N_127);
    
    \Cel_ongoing_RNO[13]\ : XA1
      port map(A => \Cel_ongoing[13]_net_1\, B => N_28_0, C => 
        N_371, Y => \Cel_ongoing_RNO[13]_net_1\);
    
    \Cel_ongoing_RNO[24]\ : NOR2A
      port map(A => N_371, B => N_63, Y => N_443);
    
    \Chanel_ongoing_RNO[16]\ : XA1C
      port map(A => \Chanel_ongoing[16]_net_1\, B => N_272, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => N_232);
    
    \Chanel_ongoing_RNI0M7B[19]\ : OR2A
      port map(A => \Chanel_ongoing[19]_net_1\, B => N_276, Y => 
        N_278);
    
    \Cel_ongoing_RNO[20]\ : NOR2A
      port map(A => N_371_0, B => N_55, Y => N_439);
    
    \Cel_ongoing[5]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[5]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[5]_net_1\);
    
    \Cel_ongoing[29]\ : DFN1C0
      port map(D => N_448, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[29]_net_1\);
    
    \IIR_CEL_STATE_i_RNIBA69[9]\ : AO1D
      port map(A => sample_val_delay, B => 
        \IIR_CEL_STATE_i[9]_net_1\, C => N_294, Y => 
        un1_IIR_CEL_STATE_20);
    
    \Chanel_ongoing_RNO_0[1]\ : XNOR2
      port map(A => \Chanel_ongoing[0]_net_1\, B => 
        \Chanel_ongoing[1]_net_1\, Y => Chanel_ongoing_n1_0_i_0_0);
    
    \Chanel_ongoing_RNO[27]\ : XA1C
      port map(A => \Chanel_ongoing[27]_net_1\, B => N_292, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n27);
    
    \waddr_previous_RNO[0]\ : OR2A
      port map(A => N_248, B => N_334, Y => un1_IIR_CEL_STATE_25);
    
    un1_IIR_CEL_STATE_17_m69 : NOR2B
      port map(A => N_68, B => \Cel_ongoing[27]_net_1\, Y => N_70);
    
    \ram_sel_Wdata[0]\ : DFN1E0C0
      port map(D => N_567_i_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => \IIR_CEL_STATE[8]_net_1\, Q => ram_sel_Wdata(0));
    
    un1_IIR_CEL_STATE_17_m74 : NOR3C
      port map(A => \Cel_ongoing[29]_net_1\, B => 
        \Cel_ongoing[30]_net_1\, C => N_72, Y => N_75);
    
    \Chanel_ongoing[4]\ : DFN1E1C0
      port map(D => N_11, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[4]_net_1\);
    
    \Cel_ongoing_RNO[0]\ : OAI1
      port map(A => N_480, B => un1_IIR_CEL_STATE_20, C => 
        \Cel_ongoing_6_i_i_1[0]\, Y => N_206);
    
    \IIR_CEL_STATE_RNI9V445_0[4]\ : OR2A
      port map(A => \IIR_CEL_STATE[4]_net_1\, B => N_328, Y => 
        N_480);
    
    \Chanel_ongoing_RNO_0[31]\ : OR2A
      port map(A => \Chanel_ongoing[30]_net_1\, B => N_327, Y => 
        N_335);
    
    \Chanel_ongoing_RNI8391[13]\ : NOR2
      port map(A => \Chanel_ongoing[13]_net_1\, B => 
        \Chanel_ongoing[22]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_6);
    
    \Chanel_ongoing_RNO_0[10]\ : AX1E
      port map(A => \Chanel_ongoing[9]_net_1\, B => N_256, C => 
        \Chanel_ongoing[10]_net_1\, Y => N_373_i);
    
    \Chanel_ongoing_RNO[8]\ : NOR2
      port map(A => Chanel_ongoing_n8_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_651);
    
    \IIR_CEL_STATE_RNIJ1T5[1]\ : OR2
      port map(A => \IIR_CEL_STATE[1]_net_1\, B => 
        \IIR_CEL_STATE[0]_net_1\, Y => N_294);
    
    \Chanel_ongoing_RNO[15]\ : XA1C
      port map(A => \Chanel_ongoing[15]_net_1\, B => N_271, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => N_229);
    
    \Chanel_ongoing[7]\ : DFN1E1C0
      port map(D => N_650, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[7]_net_1\);
    
    \Cel_ongoing_RNO[8]\ : NOR2A
      port map(A => N_371_0, B => N_38, Y => 
        \Cel_ongoing_RNO[8]_net_1\);
    
    \Cel_ongoing[13]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[13]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[13]_net_1\);
    
    \Cel_ongoing[12]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[12]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[12]_net_1\);
    
    \Chanel_ongoing_RNO[22]\ : XA1C
      port map(A => \Chanel_ongoing[22]_net_1\, B => N_725, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n22);
    
    un1_IIR_CEL_STATE_17_m65 : NOR2B
      port map(A => N_64, B => \Cel_ongoing[25]_net_1\, Y => N_66);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_1 : NOR2B
      port map(A => \Cel_ongoing[16]_net_1\, B => 
        \Cel_ongoing[17]_net_1\, Y => ADD_32x32_fast_I129_un1_Y_1);
    
    \Chanel_ongoing_RNO[28]\ : XA1C
      port map(A => \Chanel_ongoing[28]_net_1\, B => N_293, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n28);
    
    \Cel_ongoing_RNO[14]\ : NOR2A
      port map(A => N_371_0, B => \un1_IIR_CEL_STATE_17_i[17]\, Y
         => \Cel_ongoing_RNO[14]_net_1\);
    
    \Cel_ongoing_RNO[1]\ : NOR2A
      port map(A => N_371, B => N_31_0, Y => 
        \Cel_ongoing_RNO[1]_net_1\);
    
    un1_IIR_CEL_STATE_17_m33 : AX1E
      port map(A => \Cel_ongoing[3]_net_1\, B => N_18_0, C => 
        \Cel_ongoing[4]_net_1\, Y => N_34_0);
    
    \Cel_ongoing_RNO[10]\ : NOR2A
      port map(A => N_371_0, B => N_40, Y => 
        \Cel_ongoing_RNO[10]_net_1\);
    
    \Cel_ongoing_RNICE615[2]\ : OR2B
      port map(A => N_325_i, B => \Cel_ongoing[2]_net_1\, Y => 
        N_328);
    
    un1_IIR_CEL_STATE_17_m59 : NOR3C
      port map(A => \Cel_ongoing[21]_net_1\, B => N_56, C => 
        \Cel_ongoing[22]_net_1\, Y => N_60);
    
    \Chanel_ongoing_RNI7JI2[27]\ : NOR3A
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_10, B => 
        \Chanel_ongoing[28]_net_1\, C => 
        \Chanel_ongoing[27]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_20);
    
    \IIR_CEL_STATE_i_RNIDS23[9]\ : NOR2A
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, B => 
        \IIR_CEL_STATE[4]_net_1\, Y => N_733_1);
    
    \Chanel_ongoing_RNI5255[23]\ : NOR3C
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_8, B => 
        Cel_ongoing_0_sqmuxa_0_a2_0_7, C => 
        Cel_ongoing_0_sqmuxa_0_a2_0_20, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_25);
    
    \Cel_ongoing_RNIL5C8[16]\ : NOR2
      port map(A => \Cel_ongoing[15]_net_1\, B => 
        \Cel_ongoing[16]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_8[1]\);
    
    \Cel_ongoing[6]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[6]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[6]_net_1\);
    
    \IIR_CEL_STATE[3]\ : DFN1E1
      port map(D => \IIR_CEL_STATE[7]_net_1\, CLK => HCLK_c, E
         => HRESETn_c, Q => \IIR_CEL_STATE[3]_net_1\);
    
    \Cel_ongoing_RNO[29]\ : XA1
      port map(A => \Cel_ongoing[29]_net_1\, B => N_72, C => 
        N_371, Y => N_448);
    
    raddr_add1_RNO_2 : OR2A
      port map(A => N_328, B => raddr_add1_2_i_a2_0_0, Y => N_736);
    
    \Chanel_ongoing_RNI9V81[14]\ : NOR2
      port map(A => \Chanel_ongoing[14]_net_1\, B => 
        \Chanel_ongoing[15]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_11);
    
    \Chanel_ongoing[0]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[0]_net_1\);
    
    \Cel_ongoing_RNO[6]\ : NOR2A
      port map(A => N_371_0, B => N_36_0, Y => 
        \Cel_ongoing_RNO[6]_net_1\);
    
    \Cel_ongoing[14]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[14]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[14]_net_1\);
    
    \alu_selected_coeff_0_RNI679D[2]\ : XNOR2
      port map(A => S(8), B => \alu_sel_coeff_0[2]\, Y => 
        alu_selected_coeff_n2_0_i_0);
    
    un1_IIR_CEL_STATE_17_m55 : NOR3C
      port map(A => \Cel_ongoing[19]_net_1\, B => N_52, C => 
        \Cel_ongoing[20]_net_1\, Y => N_56);
    
    \Cel_ongoing[9]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[9]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[9]_net_1\);
    
    sample_in_rot : DFN1E0C0
      port map(D => sample_in_rot_2, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_353, Q => sample_in_rotate);
    
    \Chanel_ongoing_RNO[17]\ : XA1C
      port map(A => \Chanel_ongoing[17]_net_1\, B => N_273, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n17);
    
    \alu_selected_coeff[1]\ : DFN1E1C0
      port map(D => N_712, CLK => HCLK_c, CLR => HRESETn_c, E => 
        alu_selected_coeffe, Q => alu_sel_coeff(1));
    
    \Cel_ongoing[8]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[8]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[8]_net_1\);
    
    un1_IIR_CEL_STATE_17_m32 : XNOR2
      port map(A => N_18_0, B => \Cel_ongoing[3]_net_1\, Y => 
        N_33_0);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I174_Y_0 : AX1E
      port map(A => \Cel_ongoing[13]_net_1\, B => N_28_0, C => 
        \Cel_ongoing[14]_net_1\, Y => 
        \un1_IIR_CEL_STATE_17_i[17]\);
    
    \IIR_CEL_STATE[8]\ : DFN1E1
      port map(D => N_274, CLK => HCLK_c, E => HRESETn_c, Q => 
        \IIR_CEL_STATE[8]_net_1\);
    
    un1_IIR_CEL_STATE_17_m41 : AX1E
      port map(A => \Cel_ongoing[11]_net_1\, B => N_26_0, C => 
        \Cel_ongoing[12]_net_1\, Y => N_42);
    
    \raddr_add1\ : DFN1C0
      port map(D => N_723_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => raddr_add1);
    
    \IIR_CEL_STATE[1]\ : DFN1E1
      port map(D => \IIR_CEL_STATE_ns[8]\, CLK => HCLK_c, E => 
        HRESETn_c, Q => \IIR_CEL_STATE[1]_net_1\);
    
    \alu_sel_input\ : DFN1E0C0
      port map(D => alu_sel_input_1, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_IIR_CEL_STATE_20, Q => alu_sel_input);
    
    un1_IIR_CEL_STATE_17_m58 : AX1E
      port map(A => \Cel_ongoing[21]_net_1\, B => N_56, C => 
        \Cel_ongoing[22]_net_1\, Y => N_59);
    
    \ram_write\ : DFN1E0C0
      port map(D => ram_write_2, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \IIR_CEL_STATE[8]_net_1\, Q => ram_write_net_1);
    
    \IIR_CEL_STATE_i_RNO_0[9]\ : AO1D
      port map(A => sample_val_delay, B => 
        \IIR_CEL_STATE_i[9]_net_1\, C => \IIR_CEL_STATE[0]_net_1\, 
        Y => N_180);
    
    \Chanel_ongoing[10]\ : DFN1E1C0
      port map(D => N_461, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127_0, Q => \Chanel_ongoing[10]_net_1\);
    
    \in_sel_src[1]\ : DFN1E0C0
      port map(D => N_269, CLK => HCLK_c, CLR => HRESETn_c, E => 
        un1_IIR_CEL_STATE_27, Q => in_sel_src(1));
    
    \IIR_CEL_STATE_RNI9T4D5_0[4]\ : OR2A
      port map(A => N_248, B => N_566, Y => N_371);
    
    \Chanel_ongoing[17]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n17, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127_0, Q => \Chanel_ongoing[17]_net_1\);
    
    \Cel_ongoing[7]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[7]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[7]_net_1\);
    
    \Cel_ongoing_RNO[30]\ : XA1
      port map(A => \Cel_ongoing[30]_net_1\, B => I129_un1_Y, C
         => N_371, Y => N_449);
    
    \Cel_ongoing[28]\ : DFN1C0
      port map(D => N_447, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[28]_net_1\);
    
    un1_IIR_CEL_STATE_17_m39 : AX1E
      port map(A => \Cel_ongoing[9]_net_1\, B => N_24_0, C => 
        \Cel_ongoing[10]_net_1\, Y => N_40);
    
    \Chanel_ongoing_RNO[12]\ : NOR2
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0_0, B => 
        N_216_tz, Y => N_216);
    
    \Chanel_ongoing[25]\ : DFN1E1C0
      port map(D => Chanel_ongoing_n25, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_127, Q => \Chanel_ongoing[25]_net_1\);
    
    \Cel_ongoing_RNO[19]\ : XA1
      port map(A => \Cel_ongoing[19]_net_1\, B => N_52, C => 
        N_371_0, Y => N_438);
    
    \Chanel_ongoing_RNIOAVI[6]\ : OR3C
      port map(A => Cel_ongoing_0_sqmuxa_0_a2_0_26, B => 
        Cel_ongoing_0_sqmuxa_0_a2_0_25, C => 
        Cel_ongoing_0_sqmuxa_0_a2_0_27, Y => N_796_i);
    
    \Cel_ongoing_RNO[28]\ : XA1
      port map(A => \Cel_ongoing[28]_net_1\, B => N_70, C => 
        N_371, Y => N_447);
    
    \Chanel_ongoing_RNO[18]\ : XA1B
      port map(A => \Chanel_ongoing[18]_net_1\, B => N_275, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => 
        Chanel_ongoing_n18);
    
    \Cel_ongoing_RNIFEQD[4]\ : NOR2
      port map(A => \Cel_ongoing[3]_net_1\, B => 
        \Cel_ongoing[4]_net_1\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_1[1]\);
    
    \Cel_ongoing_RNIVS741[16]\ : NOR3C
      port map(A => \in_sel_src_8_i_a2_0_o2_0_8[1]\, B => 
        \in_sel_src_8_i_a2_0_o2_0_7[1]\, C => 
        \in_sel_src_8_i_a2_0_o2_0_20[1]\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_25[1]\);
    
    \Chanel_ongoing_RNO[1]\ : NOR2
      port map(A => Chanel_ongoing_n1_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_18);
    
    \Cel_ongoing[26]\ : DFN1C0
      port map(D => N_445, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[26]_net_1\);
    
    \Cel_ongoing_RNIIROG[25]\ : NOR3A
      port map(A => \in_sel_src_8_i_a2_0_o2_0_14[1]\, B => 
        \Cel_ongoing[26]_net_1\, C => \Cel_ongoing[25]_net_1\, Y
         => \in_sel_src_8_i_a2_0_o2_0_22[1]\);
    
    sample_in_rot_RNI6EV7_0 : CLKINT
      port map(A => \sample_in_rot_RNI6EV7\, Y => 
        un1_sample_in_rotate);
    
    \Chanel_ongoing[9]\ : DFN1E1C0
      port map(D => N_460, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[9]_net_1\);
    
    un1_IIR_CEL_STATE_17_m35 : AX1E
      port map(A => \Cel_ongoing[5]_net_1\, B => N_20_0, C => 
        \Cel_ongoing[6]_net_1\, Y => N_36_0);
    
    \IIR_CEL_STATE_RNIS1T5[2]\ : OR2
      port map(A => \IIR_CEL_STATE[8]_net_1\, B => 
        \IIR_CEL_STATE[2]_net_1\, Y => N_353);
    
    \Chanel_ongoing_RNO[3]\ : AO1A
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0, B => 
        N_336_i_i_0, C => \IIR_CEL_STATE_ns[8]\, Y => N_221);
    
    \Chanel_ongoing_RNO[5]\ : NOR2
      port map(A => Chanel_ongoing_n5_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_20);
    
    \Cel_ongoing_RNIJJHK2[12]\ : NOR3C
      port map(A => \in_sel_src_8_i_a2_0_o2_0_18[1]\, B => 
        \in_sel_src_8_i_a2_0_o2_0_17[1]\, C => 
        \in_sel_src_8_i_a2_0_o2_0_23[1]\, Y => 
        \in_sel_src_8_i_a2_0_o2_0_27[1]\);
    
    \alu_ctrl_RNO[1]\ : OR2
      port map(A => \IIR_CEL_STATE[8]_net_1\, B => 
        \IIR_CEL_STATE[4]_net_1\, Y => N_569);
    
    \Cel_ongoing[3]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[3]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[3]_net_1\);
    
    \Chanel_ongoing_RNO_0[2]\ : AX1C
      port map(A => \Chanel_ongoing[0]_net_1\, B => 
        \Chanel_ongoing[1]_net_1\, C => \Chanel_ongoing[2]_net_1\, 
        Y => Chanel_ongoing_n2_0_i_0_0);
    
    \Chanel_ongoing_RNO[9]\ : NOR2
      port map(A => un1_alu_sel_input_0_sqmuxa_2_i_0, B => 
        N_372_i, Y => N_460);
    
    \Cel_ongoing_RNO[18]\ : NOR2A
      port map(A => N_371_0, B => N_51, Y => N_437);
    
    \IIR_CEL_STATE[0]\ : DFN1E1
      port map(D => \IIR_CEL_STATE[1]_net_1\, CLK => HCLK_c, E
         => HRESETn_c, Q => \IIR_CEL_STATE[0]_net_1\);
    
    \Cel_ongoing[27]\ : DFN1C0
      port map(D => N_446, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[27]_net_1\);
    
    \alu_selected_coeff[2]\ : DFN1E1C0
      port map(D => N_713, CLK => HCLK_c, CLR => HRESETn_c, E => 
        alu_selected_coeffe, Q => \alu_sel_coeff[2]\);
    
    \alu_ctrl_RNO[2]\ : INV
      port map(A => \IIR_CEL_STATE_i[9]_net_1\, Y => 
        \IIR_CEL_STATE_i_i[9]\);
    
    un1_IIR_CEL_STATE_17_ADD_32x32_fast_I129_un1_Y_3 : NOR2B
      port map(A => \Cel_ongoing[20]_net_1\, B => 
        \Cel_ongoing[21]_net_1\, Y => ADD_32x32_fast_I129_un1_Y_3);
    
    \Cel_ongoing[21]\ : DFN1C0
      port map(D => N_440, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[21]_net_1\);
    
    \Chanel_ongoing_RNIBRLH[29]\ : OR2A
      port map(A => \Chanel_ongoing[29]_net_1\, B => N_295, Y => 
        N_327);
    
    sample_in_rot_RNI6EV7 : OR2
      port map(A => sample_val_delay, B => sample_in_rotate, Y
         => \sample_in_rot_RNI6EV7\);
    
    \Cel_ongoing_RNO_2[0]\ : AOI1B
      port map(A => \un1_IIR_CEL_STATE_17_i_1_i_0[31]\, B => N_6, 
        C => N_457, Y => \Cel_ongoing_6_i_i_0[0]\);
    
    \Cel_ongoing_RNO[27]\ : XA1
      port map(A => \Cel_ongoing[27]_net_1\, B => N_68, C => 
        N_371, Y => N_446);
    
    \Cel_ongoing[20]\ : DFN1C0
      port map(D => N_439, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \Cel_ongoing[20]_net_1\);
    
    \Chanel_ongoing_RNID718[14]\ : OR2A
      port map(A => \Chanel_ongoing[14]_net_1\, B => N_270, Y => 
        N_271);
    
    un1_IIR_CEL_STATE_17_m43 : NOR3C
      port map(A => \Cel_ongoing[13]_net_1\, B => N_28_0, C => 
        \Cel_ongoing[14]_net_1\, Y => N_44);
    
    \Chanel_ongoing_RNO_0[8]\ : AX1E
      port map(A => \Chanel_ongoing[7]_net_1\, B => N_254, C => 
        \Chanel_ongoing[8]_net_1\, Y => Chanel_ongoing_n8_0_i_0_0);
    
    \Cel_ongoing[1]\ : DFN1C0
      port map(D => \Cel_ongoing_RNO[1]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \Cel_ongoing[1]_net_1\);
    
    \Chanel_ongoing_RNIDV81[16]\ : NOR2
      port map(A => \Chanel_ongoing[16]_net_1\, B => 
        \Chanel_ongoing[17]_net_1\, Y => 
        Cel_ongoing_0_sqmuxa_0_a2_0_12);
    
    \Cel_ongoing_RNO[26]\ : XA1
      port map(A => \Cel_ongoing[26]_net_1\, B => N_66, C => 
        N_371, Y => N_445);
    
    \Chanel_ongoing_RNO_0[4]\ : AX1A
      port map(A => N_250, B => \Chanel_ongoing[3]_net_1\, C => 
        \Chanel_ongoing[4]_net_1\, Y => Chanel_ongoing_n4_0_i_0_0);
    
    \Chanel_ongoing_RNO[7]\ : NOR2A
      port map(A => Chanel_ongoing_n7_0_i_0_0, B => 
        un1_alu_sel_input_0_sqmuxa_2_i_0_0, Y => N_650);
    
    \waddr_previous_RNO[1]\ : OR2
      port map(A => un1_IIR_CEL_STATE_22, B => N_567_i_0, Y => 
        N_729);
    
    un1_IIR_CEL_STATE_17_m27 : NOR3C
      port map(A => \Cel_ongoing[11]_net_1\, B => N_26_0, C => 
        \Cel_ongoing[12]_net_1\, Y => N_28_0);
    
    \Chanel_ongoing_RNIFV81[17]\ : NOR2B
      port map(A => \Chanel_ongoing[17]_net_1\, B => 
        \Chanel_ongoing[18]_net_1\, Y => 
        Chanel_ongoing_n23_0_0_0_o2_m6_0_a2_2);
    
    \alu_ctrl_RNO[0]\ : OR3
      port map(A => \IIR_CEL_STATE[3]_net_1\, B => 
        \IIR_CEL_STATE[6]_net_1\, C => N_289, Y => N_568_i_0);
    
    \Chanel_ongoing_RNO[23]\ : XA1C
      port map(A => \Chanel_ongoing[23]_net_1\, B => 
        \Chanel_ongoing_RNISG5D[13]_net_1\, C => 
        un1_alu_sel_input_0_sqmuxa_2_i_0, Y => Chanel_ongoing_n23);
    
    \Chanel_ongoing[5]\ : DFN1E1C0
      port map(D => N_20, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_127, Q => \Chanel_ongoing[5]_net_1\);
    
    \Cel_ongoing_RNO_3[0]\ : OR3A
      port map(A => N_274, B => N_294, C => 
        \IIR_CEL_STATE[4]_net_1\, Y => N_457);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity IIR_CEL_CTRLR_v2 is

    port( sample_filter_v2_out_0   : out   std_logic;
          sample_filter_v2_out_1   : out   std_logic;
          sample_filter_v2_out_2   : out   std_logic;
          sample_filter_v2_out_3   : out   std_logic;
          sample_filter_v2_out_4   : out   std_logic;
          sample_filter_v2_out_5   : out   std_logic;
          sample_filter_v2_out_6   : out   std_logic;
          sample_filter_v2_out_7   : out   std_logic;
          sample_filter_v2_out_8   : out   std_logic;
          sample_filter_v2_out_9   : out   std_logic;
          sample_filter_v2_out_10  : out   std_logic;
          sample_filter_v2_out_11  : out   std_logic;
          sample_filter_v2_out_12  : out   std_logic;
          sample_filter_v2_out_13  : out   std_logic;
          sample_filter_v2_out_14  : out   std_logic;
          sample_filter_v2_out_15  : out   std_logic;
          sample_filter_v2_out_18  : out   std_logic;
          sample_filter_v2_out_19  : out   std_logic;
          sample_filter_v2_out_20  : out   std_logic;
          sample_filter_v2_out_21  : out   std_logic;
          sample_filter_v2_out_22  : out   std_logic;
          sample_filter_v2_out_23  : out   std_logic;
          sample_filter_v2_out_24  : out   std_logic;
          sample_filter_v2_out_25  : out   std_logic;
          sample_filter_v2_out_26  : out   std_logic;
          sample_filter_v2_out_27  : out   std_logic;
          sample_filter_v2_out_28  : out   std_logic;
          sample_filter_v2_out_29  : out   std_logic;
          sample_filter_v2_out_30  : out   std_logic;
          sample_filter_v2_out_31  : out   std_logic;
          sample_filter_v2_out_32  : out   std_logic;
          sample_filter_v2_out_33  : out   std_logic;
          sample_filter_v2_out_36  : out   std_logic;
          sample_filter_v2_out_37  : out   std_logic;
          sample_filter_v2_out_38  : out   std_logic;
          sample_filter_v2_out_39  : out   std_logic;
          sample_filter_v2_out_40  : out   std_logic;
          sample_filter_v2_out_41  : out   std_logic;
          sample_filter_v2_out_42  : out   std_logic;
          sample_filter_v2_out_43  : out   std_logic;
          sample_filter_v2_out_44  : out   std_logic;
          sample_filter_v2_out_45  : out   std_logic;
          sample_filter_v2_out_46  : out   std_logic;
          sample_filter_v2_out_47  : out   std_logic;
          sample_filter_v2_out_48  : out   std_logic;
          sample_filter_v2_out_49  : out   std_logic;
          sample_filter_v2_out_50  : out   std_logic;
          sample_filter_v2_out_51  : out   std_logic;
          sample_filter_v2_out_54  : out   std_logic;
          sample_filter_v2_out_55  : out   std_logic;
          sample_filter_v2_out_56  : out   std_logic;
          sample_filter_v2_out_57  : out   std_logic;
          sample_filter_v2_out_58  : out   std_logic;
          sample_filter_v2_out_59  : out   std_logic;
          sample_filter_v2_out_60  : out   std_logic;
          sample_filter_v2_out_61  : out   std_logic;
          sample_filter_v2_out_62  : out   std_logic;
          sample_filter_v2_out_63  : out   std_logic;
          sample_filter_v2_out_64  : out   std_logic;
          sample_filter_v2_out_65  : out   std_logic;
          sample_filter_v2_out_66  : out   std_logic;
          sample_filter_v2_out_67  : out   std_logic;
          sample_filter_v2_out_68  : out   std_logic;
          sample_filter_v2_out_69  : out   std_logic;
          sample_filter_v2_out_90  : out   std_logic;
          sample_filter_v2_out_91  : out   std_logic;
          sample_filter_v2_out_92  : out   std_logic;
          sample_filter_v2_out_93  : out   std_logic;
          sample_filter_v2_out_94  : out   std_logic;
          sample_filter_v2_out_95  : out   std_logic;
          sample_filter_v2_out_96  : out   std_logic;
          sample_filter_v2_out_97  : out   std_logic;
          sample_filter_v2_out_98  : out   std_logic;
          sample_filter_v2_out_99  : out   std_logic;
          sample_filter_v2_out_100 : out   std_logic;
          sample_filter_v2_out_101 : out   std_logic;
          sample_filter_v2_out_102 : out   std_logic;
          sample_filter_v2_out_103 : out   std_logic;
          sample_filter_v2_out_104 : out   std_logic;
          sample_filter_v2_out_105 : out   std_logic;
          sample_filter_v2_out_108 : out   std_logic;
          sample_filter_v2_out_126 : out   std_logic;
          sample_filter_v2_out_109 : out   std_logic;
          sample_filter_v2_out_127 : out   std_logic;
          sample_filter_v2_out_110 : out   std_logic;
          sample_filter_v2_out_128 : out   std_logic;
          sample_filter_v2_out_111 : out   std_logic;
          sample_filter_v2_out_129 : out   std_logic;
          sample_filter_v2_out_112 : out   std_logic;
          sample_filter_v2_out_130 : out   std_logic;
          sample_filter_v2_out_113 : out   std_logic;
          sample_filter_v2_out_131 : out   std_logic;
          sample_filter_v2_out_114 : out   std_logic;
          sample_filter_v2_out_132 : out   std_logic;
          sample_filter_v2_out_115 : out   std_logic;
          sample_filter_v2_out_133 : out   std_logic;
          sample_filter_v2_out_116 : out   std_logic;
          sample_filter_v2_out_134 : out   std_logic;
          sample_filter_v2_out_117 : out   std_logic;
          sample_filter_v2_out_135 : out   std_logic;
          sample_filter_v2_out_118 : out   std_logic;
          sample_filter_v2_out_136 : out   std_logic;
          sample_filter_v2_out_119 : out   std_logic;
          sample_filter_v2_out_137 : out   std_logic;
          sample_filter_v2_out_120 : out   std_logic;
          sample_filter_v2_out_138 : out   std_logic;
          sample_filter_v2_out_121 : out   std_logic;
          sample_filter_v2_out_139 : out   std_logic;
          sample_filter_v2_out_122 : out   std_logic;
          sample_filter_v2_out_140 : out   std_logic;
          sample_filter_v2_out_123 : out   std_logic;
          sample_filter_v2_out_141 : out   std_logic;
          sample_6                 : in    std_logic_vector(15 downto 0);
          sample_5                 : in    std_logic_vector(15 downto 0);
          sample_2                 : in    std_logic_vector(15 downto 0);
          sample_0                 : in    std_logic_vector(15 downto 0);
          sample_1                 : in    std_logic_vector(15 downto 0);
          sample_3                 : in    std_logic_vector(15 downto 0);
          sample_4                 : in    std_logic_vector(15 downto 0);
          sample_7                 : in    std_logic_vector(15 downto 0);
          IIR_CEL_CTRLR_v2_VCC     : in    std_logic;
          IIR_CEL_CTRLR_v2_GND     : in    std_logic;
          HRESETn_c                : in    std_logic;
          HCLK_c                   : in    std_logic;
          sample_filter_v2_out_val : out   std_logic;
          sample_val_delay         : in    std_logic
        );

end IIR_CEL_CTRLR_v2;

architecture DEF_ARCH of IIR_CEL_CTRLR_v2 is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component IIR_CEL_CTRLR_v2_DATAFLOW
    port( alu_ctrl                      : in    std_logic_vector(2 downto 0) := (others => 'U');
          S                             : out   std_logic_vector(8 to 8);
          S_i_0                         : out   std_logic_vector(33 to 33);
          alu_sel_coeff                 : in    std_logic_vector(4 downto 0) := (others => 'U');
          alu_sel_coeff_0_2             : in    std_logic := 'U';
          alu_sel_coeff_0_0             : in    std_logic := 'U';
          waddr_previous                : in    std_logic_vector(1 downto 0) := (others => 'U');
          sample_0                      : in    std_logic_vector(14 downto 0) := (others => 'U');
          sample_in_buf                 : in    std_logic_vector(143 downto 129) := (others => 'U');
          ram_sel_Wdata                 : in    std_logic_vector(1 downto 0) := (others => 'U');
          sample_out_s_0                : out   std_logic;
          sample_out_s_1                : out   std_logic;
          sample_out_s_3                : out   std_logic;
          sample_out_s_2                : out   std_logic;
          sample_out_s_10               : out   std_logic;
          sample_out_s_15               : out   std_logic;
          sample_out_s_14               : out   std_logic;
          sample_out_s_13               : out   std_logic;
          sample_out_s_12               : out   std_logic;
          sample_out_s_11               : out   std_logic;
          sample_out_s_9                : out   std_logic;
          sample_out_s_8                : out   std_logic;
          sample_out_s_7                : out   std_logic;
          sample_out_s_6                : out   std_logic;
          sample_out_s_5                : out   std_logic;
          sample_out_s_4                : out   std_logic;
          sample_in_s_1                 : in    std_logic_vector(17 to 17) := (others => 'U');
          in_sel_src                    : in    std_logic_vector(1 downto 0) := (others => 'U');
          raddr_rst                     : in    std_logic := 'U';
          raddr_add1                    : in    std_logic := 'U';
          ram_write                     : in    std_logic := 'U';
          IIR_CEL_CTRLR_v2_DATAFLOW_GND : in    std_logic := 'U';
          IIR_CEL_CTRLR_v2_DATAFLOW_VCC : in    std_logic := 'U';
          ram_write_i                   : in    std_logic := 'U';
          HRESETn_c                     : in    std_logic := 'U';
          HCLK_c                        : in    std_logic := 'U';
          sample_val_delay              : in    std_logic := 'U';
          alu_sel_input                 : in    std_logic := 'U'
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component IIR_CEL_CTRLR_v2_CONTROL
    port( alu_ctrl             : out   std_logic_vector(2 downto 0);
          ram_sel_Wdata        : out   std_logic_vector(1 downto 0);
          waddr_previous       : out   std_logic_vector(1 downto 0);
          in_sel_src           : out   std_logic_vector(1 downto 0);
          S_i_0                : in    std_logic_vector(33 to 33) := (others => 'U');
          S                    : in    std_logic_vector(8 to 8) := (others => 'U');
          alu_sel_coeff        : out   std_logic_vector(4 downto 0);
          alu_sel_coeff_0_2    : out   std_logic;
          alu_sel_coeff_0_0    : out   std_logic;
          sample_out_rot_s     : out   std_logic;
          sample_out_val_s     : out   std_logic;
          raddr_rst            : out   std_logic;
          alu_sel_input        : out   std_logic;
          raddr_add1           : out   std_logic;
          sample_val_delay     : in    std_logic := 'U';
          ram_write            : out   std_logic;
          ram_write_i          : out   std_logic;
          un1_sample_in_rotate : out   std_logic;
          sample_out_rot_s_0   : out   std_logic;
          sample_out_rot_s_1   : out   std_logic;
          sample_out_rot_s_2   : out   std_logic;
          sample_out_rot_s_3   : out   std_logic;
          sample_out_rot_s_4   : out   std_logic;
          HRESETn_c            : in    std_logic := 'U';
          HCLK_c               : in    std_logic := 'U'
        );
  end component;

    signal \sample_in_buf_581[9]\, \sample_in_buf[135]\, 
        \sample_in_buf_349[59]\, \sample_in_buf[41]\, 
        \sample_in_buf_669[64]\, \sample_in_buf[46]\, 
        \sample_in_buf_293[76]\, \sample_in_buf[58]\, 
        \sample_in_buf_501[115]\, \sample_in_buf[97]\, 
        \sample_in_buf_821[120]\, \sample_in_buf[102]\, 
        \sample_in_buf_637[135]\, \sample_in_buf[117]\, 
        \sample_in_buf_965[15]\, \sample_in_buf[141]\, 
        \sample_in_buf_29[54]\, \sample_in_buf[36]\, 
        \sample_in_buf_285[58]\, \sample_in_buf[40]\, 
        \sample_in_buf_813[102]\, \sample_in_buf[84]\, 
        \sample_in_buf_437[114]\, \sample_in_buf[96]\, 
        \sample_in_buf_1021[141]\, \sample_in_buf[123]\, 
        \sample_in_buf_645[10]\, \sample_in_buf[136]\, 
        \sample_in_buf_853[49]\, \sample_in_buf[31]\, 
        \sample_in_buf_1045[52]\, \sample_in_buf[34]\, 
        \sample_in_buf_805[84]\, \sample_in_buf[66]\, 
        \sample_in_buf_493[97]\, \sample_in_buf[79]\, 
        \sample_in_buf_701[136]\, \sample_in_buf[118]\, 
        \sample_in_buf_389[6]\, \sample_in_buf[132]\, 
        \sample_in_buf_341[41]\, \sample_in_buf[23]\, 
        \sample_in_buf_605[63]\, \sample_in_buf[45]\, 
        \sample_in_buf_1117[71]\, \sample_in_buf[53]\, 
        \sample_in_buf_757[119]\, \sample_in_buf[101]\, 
        \sample_in_buf_445[132]\, \sample_in_buf[114]\, 
        \sample_in_buf_277[40]\, \sample_in_buf[22]\, 
        \sample_in_buf_725[47]\, \sample_in_buf[29]\, 
        \sample_in_buf_421[78]\, \sample_in_buf[60]\, 
        \sample_in_buf_373[113]\, \sample_in_buf[95]\, 
        \sample_in_buf_1013[123]\, \sample_in_buf[105]\, 
        \sample_in_buf_261[4]\, \sample_in_buf[130]\, 
        \sample_in_buf_21[36]\, \sample_in_buf[18]\, 
        \sample_in_buf_221[57]\, \sample_in_buf[39]\, 
        \sample_in_buf_749[101]\, \sample_in_buf[83]\, 
        \sample_in_buf_1133[107]\, \sample_in_buf[89]\, 
        \sample_in_buf_317[130]\, \sample_in_buf[112]\, 
        \sample_in_buf_517[8]\, \sample_in_buf[134]\, 
        \sample_in_buf_773[12]\, \sample_in_buf[138]\, 
        \sample_in_buf_1101[35]\, \sample_in_buf[17]\, 
        \sample_in_buf_213[39]\, \sample_in_buf[21]\, 
        \sample_in_buf_477[61]\, \sample_in_buf[43]\, 
        \sample_in_buf_1069[106]\, \sample_in_buf[88]\, 
        \sample_in_buf_573[134]\, \sample_in_buf[116]\, 
        \sample_in_buf_829[138]\, \sample_in_buf[120]\, 
        \sample_in_buf_325[5]\, \sample_in_buf[131]\, 
        \sample_in_buf_845[31]\, \sample_in_buf[13]\, 
        \sample_in_buf_909[32]\, \sample_in_buf[14]\, 
        \sample_in_buf_981[51]\, \sample_in_buf[33]\, 
        \sample_in_buf_741[83]\, \sample_in_buf[65]\, 
        \sample_in_buf_933[86]\, \sample_in_buf[68]\, 
        \sample_in_buf_1125[89]\, \sample_in_buf[71]\, 
        \sample_in_buf_237[93]\, \sample_in_buf[75]\, 
        \sample_in_buf_245[111]\, \sample_in_buf[93]\, 
        \sample_in_buf_381[131]\, \sample_in_buf[113]\, 
        \sample_in_buf_781[30]\, \sample_in_buf[12]\, 
        \sample_in_buf_789[48]\, \sample_in_buf[30]\, 
        \sample_in_buf_917[50]\, \sample_in_buf[32]\, 
        \sample_in_buf_549[80]\, \sample_in_buf[62]\, 
        \sample_in_buf_613[81]\, \sample_in_buf[63]\, 
        \sample_in_buf_997[87]\, \sample_in_buf[69]\, 
        \sample_in_buf_365[95]\, \sample_in_buf[77]\, 
        \sample_in_buf_949[122]\, \sample_in_buf[104]\, 
        \sample_in_buf_837[13]\, \sample_in_buf[139]\, 
        \sample_in_buf_653[28]\, \sample_in_buf[10]\, 
        \sample_in_buf_469[43]\, \sample_in_buf[25]\, 
        \sample_in_buf_37[72]\, \sample_in_buf[54]\, 
        \sample_in_buf_877[103]\, \sample_in_buf[85]\, 
        \sample_in_buf_893[139]\, \sample_in_buf[121]\, 
        \sample_in_buf_589[27]\, \sample_in_buf[9]\, 
        \sample_in_buf_973[33]\, \sample_in_buf[15]\, 
        \sample_in_buf_533[44]\, \sample_in_buf[26]\, 
        \sample_in_buf_861[67]\, \sample_in_buf[49]\, 
        \sample_in_buf_989[69]\, \sample_in_buf[51]\, 
        \sample_in_buf_869[85]\, \sample_in_buf[67]\, 
        \sample_in_buf_45[90]\, \sample_in_buf[72]\, 
        \sample_in_buf_301[94]\, \sample_in_buf[76]\, 
        \sample_in_buf_941[104]\, \sample_in_buf[86]\, 
        \sample_in_buf_565[116]\, \sample_in_buf[98]\, 
        \sample_in_buf_197[3]\, \sample_in_buf[129]\, 
        \sample_in_buf_525[26]\, \sample_in_buf[8]\, 
        \sample_in_buf_405[42]\, \sample_in_buf[24]\, 
        \sample_in_buf_797[66]\, \sample_in_buf[48]\, 
        \sample_in_buf_677[82]\, \sample_in_buf[64]\, 
        \sample_in_buf_1141[125]\, \sample_in_buf[107]\, 
        \sample_in_buf_253[129]\, \sample_in_buf[111]\, 
        \sample_in_buf_901[14]\, \sample_in_buf[140]\, 
        \sample_in_buf_1029[16]\, \sample_in_buf[142]\, 
        \sample_in_buf_461[25]\, \sample_in_buf[7]\, 
        \sample_in_buf_1037[34]\, \sample_in_buf[16]\, 
        \sample_in_buf_429[96]\, \sample_in_buf[78]\, 
        \sample_in_buf_957[140]\, \sample_in_buf[122]\, 
        \sample_in_buf_1085[142]\, \sample_in_buf[124]\, 
        \sample_in_buf_709[11]\, \sample_in_buf[137]\, 
        \sample_in_buf_397[24]\, \sample_in_buf[6]\, 
        \sample_in_buf_733[65]\, \sample_in_buf[47]\, 
        \sample_in_buf_485[79]\, \sample_in_buf[61]\, 
        \sample_in_buf_1077[124]\, \sample_in_buf[106]\, 
        \sample_in_buf_765[137]\, \sample_in_buf[119]\, 
        \sample_in_buf_269[22]\, \sample_in_buf[4]\, 
        \sample_in_buf_333[23]\, \sample_in_buf[5]\, 
        \sample_in_buf_597[45]\, \sample_in_buf[27]\, 
        \sample_in_buf_541[62]\, \sample_in_buf[44]\, 
        \sample_in_buf_925[68]\, \sample_in_buf[50]\, 
        \sample_in_buf_1053[70]\, \sample_in_buf[52]\, 
        \sample_in_buf_1061[88]\, \sample_in_buf[70]\, 
        \sample_in_buf_557[98]\, \sample_in_buf[80]\, 
        \sample_in_buf_621[99]\, \sample_in_buf[81]\, 
        \sample_in_buf_309[112]\, \sample_in_buf[94]\, 
        \sample_in_buf_629[117]\, \sample_in_buf[99]\, 
        \sample_in_buf_693[118]\, \sample_in_buf[100]\, 
        \sample_in_buf_5[0]\, \sample_in_buf[128]\, 
        \sample_in_buf_205[21]\, \sample_in_buf[3]\, 
        \sample_in_buf_413[60]\, \sample_in_buf[42]\, 
        \sample_in_buf_1005[105]\, \sample_in_buf[87]\, 
        \sample_in_buf_61[126]\, \sample_in_buf[108]\, 
        \sample_in_s_1[17]\, \sample_in_buf_453[7]\, 
        \sample_in_buf[133]\, \sample_in_buf_13[18]\, 
        \sample_in_buf[0]\, \sample_in_buf_717[29]\, 
        \sample_in_buf[11]\, \sample_in_buf_661[46]\, 
        \sample_in_buf[28]\, \sample_in_buf_1109[53]\, 
        \sample_in_buf[35]\, \sample_in_buf_229[75]\, 
        \sample_in_buf[57]\, \sample_in_buf_357[77]\, 
        \sample_in_buf[59]\, \sample_in_buf_685[100]\, 
        \sample_in_buf[82]\, \sample_in_buf_53[108]\, 
        \sample_in_buf[90]\, \sample_in_buf_885[121]\, 
        \sample_in_buf[103]\, \sample_in_buf_509[133]\, 
        \sample_in_buf[115]\, \sample_in_buf_1149[143]\, 
        \sample_in_buf[125]\, \sample_in_buf_1093[17]\, 
        \sample_in_buf[143]\, \sample_out_val_s2\, 
        sample_out_val_s, sample_out_rot_s_0, sample_out_rot_s_1, 
        \sample_filter_v2_out[125]\, \sample_filter_v2_out[124]\, 
        \sample_filter_v2_out[123]\, \sample_filter_v2_out[122]\, 
        \sample_filter_v2_out[121]\, \sample_filter_v2_out[120]\, 
        \sample_filter_v2_out[119]\, sample_out_rot_s_2, 
        \sample_filter_v2_out[118]\, \sample_filter_v2_out[117]\, 
        \sample_filter_v2_out[116]\, \sample_filter_v2_out[115]\, 
        \sample_filter_v2_out[114]\, \sample_filter_v2_out[113]\, 
        \sample_filter_v2_out[112]\, \sample_filter_v2_out[111]\, 
        \sample_filter_v2_out[110]\, \sample_filter_v2_out[107]\, 
        \sample_filter_v2_out[89]\, \sample_filter_v2_out[106]\, 
        \sample_filter_v2_out[88]\, \sample_filter_v2_out[105]\, 
        \sample_filter_v2_out[87]\, \sample_filter_v2_out[104]\, 
        \sample_filter_v2_out[86]\, \sample_filter_v2_out[103]\, 
        \sample_filter_v2_out[85]\, \sample_filter_v2_out[102]\, 
        \sample_filter_v2_out[84]\, \sample_filter_v2_out[101]\, 
        \sample_filter_v2_out[83]\, \sample_filter_v2_out[100]\, 
        \sample_filter_v2_out[82]\, \sample_filter_v2_out[99]\, 
        \sample_filter_v2_out[81]\, \sample_filter_v2_out[98]\, 
        \sample_filter_v2_out[80]\, \sample_filter_v2_out[97]\, 
        \sample_filter_v2_out[79]\, \sample_filter_v2_out[96]\, 
        \sample_filter_v2_out[78]\, \sample_filter_v2_out[95]\, 
        \sample_filter_v2_out[77]\, \sample_filter_v2_out[94]\, 
        \sample_filter_v2_out[76]\, \sample_filter_v2_out[93]\, 
        \sample_filter_v2_out[75]\, \sample_filter_v2_out[92]\, 
        \sample_filter_v2_out[74]\, sample_out_rot_s_3, 
        \sample_filter_v2_out[71]\, \sample_filter_v2_out[70]\, 
        \sample_filter_v2_out[69]\, sample_out_rot_s_4, 
        \sample_filter_v2_out[68]\, \sample_filter_v2_out[67]\, 
        \sample_filter_v2_out[66]\, \sample_filter_v2_out[65]\, 
        \sample_filter_v2_out[64]\, \sample_filter_v2_out[63]\, 
        \sample_filter_v2_out[62]\, \sample_filter_v2_out[61]\, 
        \sample_filter_v2_out[60]\, \sample_filter_v2_out[59]\, 
        \sample_filter_v2_out[58]\, \sample_filter_v2_out[57]\, 
        \sample_filter_v2_out[56]\, \sample_filter_v2_out[53]\, 
        \sample_filter_v2_out[52]\, \sample_filter_v2_out[51]\, 
        \sample_filter_v2_out[50]\, \sample_filter_v2_out[49]\, 
        \sample_filter_v2_out[48]\, \sample_filter_v2_out[47]\, 
        \sample_filter_v2_out[46]\, \sample_filter_v2_out[45]\, 
        sample_out_rot_s, \sample_filter_v2_out[44]\, 
        \sample_filter_v2_out[43]\, \sample_filter_v2_out[42]\, 
        \sample_filter_v2_out[41]\, \sample_filter_v2_out[40]\, 
        \sample_filter_v2_out[39]\, \sample_filter_v2_out[38]\, 
        un1_sample_in_rotate, \sample_filter_v2_out[35]\, 
        \sample_filter_v2_out[34]\, \sample_filter_v2_out[33]\, 
        \sample_filter_v2_out[32]\, \sample_filter_v2_out[31]\, 
        \sample_filter_v2_out[30]\, \sample_filter_v2_out[29]\, 
        \sample_filter_v2_out[28]\, \sample_filter_v2_out[27]\, 
        \sample_filter_v2_out[26]\, \sample_filter_v2_out[25]\, 
        \sample_filter_v2_out[24]\, \sample_filter_v2_out[23]\, 
        \sample_filter_v2_out[22]\, \sample_filter_v2_out[21]\, 
        \sample_filter_v2_out[20]\, \sample_filter_v2_out[17]\, 
        \sample_out_s[0]\, \sample_filter_v2_out[16]\, 
        \sample_out_s[1]\, \sample_filter_v2_out[15]\, 
        \sample_out_s[2]\, \sample_filter_v2_out[14]\, 
        \sample_out_s[3]\, \sample_filter_v2_out[13]\, 
        \sample_out_s[4]\, \sample_filter_v2_out[12]\, 
        \sample_out_s[5]\, \sample_filter_v2_out[11]\, 
        \sample_out_s[6]\, \sample_filter_v2_out[10]\, 
        \sample_out_s[7]\, \sample_filter_v2_out[9]\, 
        \sample_out_s[8]\, \sample_filter_v2_out[8]\, 
        \sample_out_s[9]\, \sample_filter_v2_out[7]\, 
        \sample_out_s[10]\, \sample_filter_v2_out[6]\, 
        \sample_out_s[11]\, \sample_filter_v2_out[5]\, 
        \sample_out_s[12]\, \sample_filter_v2_out[4]\, 
        \sample_out_s[13]\, \sample_filter_v2_out[3]\, 
        \sample_out_s[14]\, \sample_filter_v2_out[2]\, 
        \sample_out_s[15]\, \alu_ctrl[0]\, \alu_ctrl[1]\, 
        \alu_ctrl[2]\, \S[8]\, \S_i_0[33]\, \alu_sel_coeff[0]\, 
        \alu_sel_coeff[1]\, \alu_sel_coeff[2]\, 
        \alu_sel_coeff[3]\, \alu_sel_coeff[4]\, 
        \alu_sel_coeff_0[2]\, \alu_sel_coeff_0[0]\, 
        \waddr_previous[0]\, \waddr_previous[1]\, 
        \ram_sel_Wdata[0]\, \ram_sel_Wdata[1]\, \in_sel_src[0]\, 
        \in_sel_src[1]\, raddr_rst, raddr_add1, ram_write, 
        ram_write_i, alu_sel_input, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : IIR_CEL_CTRLR_v2_DATAFLOW
	Use entity work.IIR_CEL_CTRLR_v2_DATAFLOW(DEF_ARCH);
    for all : IIR_CEL_CTRLR_v2_CONTROL
	Use entity work.IIR_CEL_CTRLR_v2_CONTROL(DEF_ARCH);
begin 

    sample_filter_v2_out_0 <= \sample_filter_v2_out[2]\;
    sample_filter_v2_out_1 <= \sample_filter_v2_out[3]\;
    sample_filter_v2_out_2 <= \sample_filter_v2_out[4]\;
    sample_filter_v2_out_3 <= \sample_filter_v2_out[5]\;
    sample_filter_v2_out_4 <= \sample_filter_v2_out[6]\;
    sample_filter_v2_out_5 <= \sample_filter_v2_out[7]\;
    sample_filter_v2_out_6 <= \sample_filter_v2_out[8]\;
    sample_filter_v2_out_7 <= \sample_filter_v2_out[9]\;
    sample_filter_v2_out_8 <= \sample_filter_v2_out[10]\;
    sample_filter_v2_out_9 <= \sample_filter_v2_out[11]\;
    sample_filter_v2_out_10 <= \sample_filter_v2_out[12]\;
    sample_filter_v2_out_11 <= \sample_filter_v2_out[13]\;
    sample_filter_v2_out_12 <= \sample_filter_v2_out[14]\;
    sample_filter_v2_out_13 <= \sample_filter_v2_out[15]\;
    sample_filter_v2_out_14 <= \sample_filter_v2_out[16]\;
    sample_filter_v2_out_15 <= \sample_filter_v2_out[17]\;
    sample_filter_v2_out_18 <= \sample_filter_v2_out[20]\;
    sample_filter_v2_out_19 <= \sample_filter_v2_out[21]\;
    sample_filter_v2_out_20 <= \sample_filter_v2_out[22]\;
    sample_filter_v2_out_21 <= \sample_filter_v2_out[23]\;
    sample_filter_v2_out_22 <= \sample_filter_v2_out[24]\;
    sample_filter_v2_out_23 <= \sample_filter_v2_out[25]\;
    sample_filter_v2_out_24 <= \sample_filter_v2_out[26]\;
    sample_filter_v2_out_25 <= \sample_filter_v2_out[27]\;
    sample_filter_v2_out_26 <= \sample_filter_v2_out[28]\;
    sample_filter_v2_out_27 <= \sample_filter_v2_out[29]\;
    sample_filter_v2_out_28 <= \sample_filter_v2_out[30]\;
    sample_filter_v2_out_29 <= \sample_filter_v2_out[31]\;
    sample_filter_v2_out_30 <= \sample_filter_v2_out[32]\;
    sample_filter_v2_out_31 <= \sample_filter_v2_out[33]\;
    sample_filter_v2_out_32 <= \sample_filter_v2_out[34]\;
    sample_filter_v2_out_33 <= \sample_filter_v2_out[35]\;
    sample_filter_v2_out_36 <= \sample_filter_v2_out[38]\;
    sample_filter_v2_out_37 <= \sample_filter_v2_out[39]\;
    sample_filter_v2_out_38 <= \sample_filter_v2_out[40]\;
    sample_filter_v2_out_39 <= \sample_filter_v2_out[41]\;
    sample_filter_v2_out_40 <= \sample_filter_v2_out[42]\;
    sample_filter_v2_out_41 <= \sample_filter_v2_out[43]\;
    sample_filter_v2_out_42 <= \sample_filter_v2_out[44]\;
    sample_filter_v2_out_43 <= \sample_filter_v2_out[45]\;
    sample_filter_v2_out_44 <= \sample_filter_v2_out[46]\;
    sample_filter_v2_out_45 <= \sample_filter_v2_out[47]\;
    sample_filter_v2_out_46 <= \sample_filter_v2_out[48]\;
    sample_filter_v2_out_47 <= \sample_filter_v2_out[49]\;
    sample_filter_v2_out_48 <= \sample_filter_v2_out[50]\;
    sample_filter_v2_out_49 <= \sample_filter_v2_out[51]\;
    sample_filter_v2_out_50 <= \sample_filter_v2_out[52]\;
    sample_filter_v2_out_51 <= \sample_filter_v2_out[53]\;
    sample_filter_v2_out_54 <= \sample_filter_v2_out[56]\;
    sample_filter_v2_out_55 <= \sample_filter_v2_out[57]\;
    sample_filter_v2_out_56 <= \sample_filter_v2_out[58]\;
    sample_filter_v2_out_57 <= \sample_filter_v2_out[59]\;
    sample_filter_v2_out_58 <= \sample_filter_v2_out[60]\;
    sample_filter_v2_out_59 <= \sample_filter_v2_out[61]\;
    sample_filter_v2_out_60 <= \sample_filter_v2_out[62]\;
    sample_filter_v2_out_61 <= \sample_filter_v2_out[63]\;
    sample_filter_v2_out_62 <= \sample_filter_v2_out[64]\;
    sample_filter_v2_out_63 <= \sample_filter_v2_out[65]\;
    sample_filter_v2_out_64 <= \sample_filter_v2_out[66]\;
    sample_filter_v2_out_65 <= \sample_filter_v2_out[67]\;
    sample_filter_v2_out_66 <= \sample_filter_v2_out[68]\;
    sample_filter_v2_out_67 <= \sample_filter_v2_out[69]\;
    sample_filter_v2_out_68 <= \sample_filter_v2_out[70]\;
    sample_filter_v2_out_69 <= \sample_filter_v2_out[71]\;
    sample_filter_v2_out_90 <= \sample_filter_v2_out[92]\;
    sample_filter_v2_out_91 <= \sample_filter_v2_out[93]\;
    sample_filter_v2_out_92 <= \sample_filter_v2_out[94]\;
    sample_filter_v2_out_93 <= \sample_filter_v2_out[95]\;
    sample_filter_v2_out_94 <= \sample_filter_v2_out[96]\;
    sample_filter_v2_out_95 <= \sample_filter_v2_out[97]\;
    sample_filter_v2_out_96 <= \sample_filter_v2_out[98]\;
    sample_filter_v2_out_97 <= \sample_filter_v2_out[99]\;
    sample_filter_v2_out_98 <= \sample_filter_v2_out[100]\;
    sample_filter_v2_out_99 <= \sample_filter_v2_out[101]\;
    sample_filter_v2_out_100 <= \sample_filter_v2_out[102]\;
    sample_filter_v2_out_101 <= \sample_filter_v2_out[103]\;
    sample_filter_v2_out_102 <= \sample_filter_v2_out[104]\;
    sample_filter_v2_out_103 <= \sample_filter_v2_out[105]\;
    sample_filter_v2_out_104 <= \sample_filter_v2_out[106]\;
    sample_filter_v2_out_105 <= \sample_filter_v2_out[107]\;
    sample_filter_v2_out_108 <= \sample_filter_v2_out[110]\;
    sample_filter_v2_out_109 <= \sample_filter_v2_out[111]\;
    sample_filter_v2_out_110 <= \sample_filter_v2_out[112]\;
    sample_filter_v2_out_111 <= \sample_filter_v2_out[113]\;
    sample_filter_v2_out_112 <= \sample_filter_v2_out[114]\;
    sample_filter_v2_out_113 <= \sample_filter_v2_out[115]\;
    sample_filter_v2_out_114 <= \sample_filter_v2_out[116]\;
    sample_filter_v2_out_115 <= \sample_filter_v2_out[117]\;
    sample_filter_v2_out_116 <= \sample_filter_v2_out[118]\;
    sample_filter_v2_out_117 <= \sample_filter_v2_out[119]\;
    sample_filter_v2_out_118 <= \sample_filter_v2_out[120]\;
    sample_filter_v2_out_119 <= \sample_filter_v2_out[121]\;
    sample_filter_v2_out_120 <= \sample_filter_v2_out[122]\;
    sample_filter_v2_out_121 <= \sample_filter_v2_out[123]\;
    sample_filter_v2_out_122 <= \sample_filter_v2_out[124]\;
    sample_filter_v2_out_123 <= \sample_filter_v2_out[125]\;

    \loop_all_sample.2.loop_all_chanel.6.sample_in_buf[33]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_973[33]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[33]\);
    
    \loop_all_sample.13.loop_all_chanel.7.sample_in_buf[4]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_261[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[4]\);
    
    \loop_all_sample.9.loop_all_chanel.4.sample_in_buf_RNO[62]\ : 
        MX2
      port map(A => \sample_in_buf[44]\, B => sample_4(9), S => 
        sample_val_delay, Y => \sample_in_buf_541[62]\);
    
    \loop_all_sample.10.loop_all_chanel.2.sample_in_buf_RNO[97]\ : 
        MX2
      port map(A => \sample_in_buf[79]\, B => sample_2(10), S => 
        sample_val_delay, Y => \sample_in_buf_493[97]\);
    
    \chanel_more.all_chanel.2.all_bit.3.sample_out_s2[122]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[104]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[122]\);
    
    \loop_all_sample.5.loop_all_chanel.4.sample_in_buf_RNO[66]\ : 
        MX2
      port map(A => \sample_in_buf[48]\, B => sample_4(5), S => 
        sample_val_delay, Y => \sample_in_buf_797[66]\);
    
    \loop_all_sample.1.loop_all_chanel.6.sample_in_buf[34]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1037[34]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[34]\);
    
    \chanel_more.all_chanel.3.all_bit.1.sample_out_s2[106]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[88]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[106]\);
    
    \loop_all_sample.6.loop_all_chanel.1.sample_in_buf_RNO[119]\ : 
        MX2
      port map(A => \sample_in_buf[101]\, B => sample_1(6), S => 
        sample_val_delay, Y => \sample_in_buf_757[119]\);
    
    \loop_all_sample.12.loop_all_chanel.4.sample_in_buf_RNO[59]\ : 
        MX2
      port map(A => \sample_in_buf[41]\, B => sample_4(12), S => 
        sample_val_delay, Y => \sample_in_buf_349[59]\);
    
    \chanel_more.all_chanel.1.all_bit.6.sample_out_s2[137]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[119]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_135);
    
    \chanel_more.all_chanel.7.all_bit.3.sample_out_s2[32]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[14]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[32]\);
    
    \chanel_more.all_chanel.5.all_bit.10.sample_out_s2[61]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[43]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[61]\);
    
    \loop_all_sample.6.loop_all_chanel.0.sample_in_buf_RNO[137]\ : 
        MX2
      port map(A => \sample_in_buf[119]\, B => sample_0(6), S => 
        sample_val_delay, Y => \sample_in_buf_765[137]\);
    
    \chanel_more.all_chanel.6.all_bit.0.sample_out_s2[53]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[35]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[53]\);
    
    \chanel_more.all_chanel.4.all_bit.13.sample_out_s2[76]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[58]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[76]\);
    
    \loop_all_sample.9.loop_all_chanel.0.sample_in_buf_RNO[134]\ : 
        MX2
      port map(A => \sample_in_buf[116]\, B => sample_0(9), S => 
        sample_val_delay, Y => \sample_in_buf_573[134]\);
    
    \loop_all_sample.8.loop_all_chanel.2.sample_in_buf[99]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_621[99]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[99]\);
    
    \chanel_more.all_chanel.3.all_bit.11.sample_out_s2[96]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[78]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[96]\);
    
    \chanel_more.all_chanel.6.all_bit.2.sample_out_s2[51]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[33]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[51]\);
    
    \loop_all_sample.12.loop_all_chanel.5.sample_in_buf_RNO[41]\ : 
        MX2
      port map(A => \sample_in_buf[23]\, B => sample_5(12), S => 
        sample_val_delay, Y => \sample_in_buf_341[41]\);
    
    \loop_all_sample.1.loop_all_chanel.2.sample_in_buf[106]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1069[106]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[106]\);
    
    \loop_all_sample.17.loop_all_chanel.7.sample_in_buf_RNO[0]\ : 
        MX2
      port map(A => \sample_in_buf[128]\, B => sample_7(15), S
         => sample_val_delay, Y => \sample_in_buf_5[0]\);
    
    \loop_all_sample.13.loop_all_chanel.5.sample_in_buf[40]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_277[40]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[40]\);
    
    \loop_all_sample.13.loop_all_chanel.0.sample_in_buf_RNO[130]\ : 
        MX2
      port map(A => \sample_in_buf[112]\, B => sample_0(13), S
         => sample_val_delay, Y => \sample_in_buf_317[130]\);
    
    \loop_all_sample.3.loop_all_chanel.4.sample_in_buf_RNO[68]\ : 
        MX2
      port map(A => \sample_in_buf[50]\, B => sample_4(3), S => 
        sample_val_delay, Y => \sample_in_buf_925[68]\);
    
    \chanel_more.all_chanel.1.all_bit.3.sample_out_s2[140]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[122]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_138);
    
    \loop_all_sample.13.loop_all_chanel.2.sample_in_buf_RNO[94]\ : 
        MX2
      port map(A => \sample_in_buf[76]\, B => sample_2(13), S => 
        sample_val_delay, Y => \sample_in_buf_301[94]\);
    
    \loop_all_sample.11.loop_all_chanel.3.sample_in_buf_RNO[78]\ : 
        MX2
      port map(A => \sample_in_buf[60]\, B => sample_3(11), S => 
        sample_val_delay, Y => \sample_in_buf_421[78]\);
    
    \chanel_more.all_chanel.4.all_bit.1.sample_out_s2[88]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[70]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[88]\);
    
    \chanel_more.all_chanel.3.all_bit.4.sample_out_s2[103]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[85]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[103]\);
    
    \loop_all_sample.7.loop_all_chanel.4.sample_in_buf_RNO[64]\ : 
        MX2
      port map(A => \sample_in_buf[46]\, B => sample_4(7), S => 
        sample_val_delay, Y => \sample_in_buf_669[64]\);
    
    \loop_all_sample.5.loop_all_chanel.3.sample_in_buf[84]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_805[84]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[84]\);
    
    \chanel_more.all_chanel.6.all_bit.15.sample_out_s2[38]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[20]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[38]\);
    
    \loop_all_sample.12.loop_all_chanel.5.sample_in_buf[41]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_341[41]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[41]\);
    
    \chanel_more.all_chanel.5.all_bit.7.sample_out_s2[64]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[46]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[64]\);
    
    \chanel_more.all_chanel.5.all_bit.6.sample_out_s2[65]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[47]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[65]\);
    
    \chanel_more.all_chanel.7.all_bit.2.sample_out_s2[33]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[15]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[33]\);
    
    \loop_all_sample.9.loop_all_chanel.3.sample_in_buf_RNO[80]\ : 
        MX2
      port map(A => \sample_in_buf[62]\, B => sample_3(9), S => 
        sample_val_delay, Y => \sample_in_buf_549[80]\);
    
    \loop_all_sample.2.loop_all_chanel.4.sample_in_buf_RNO[69]\ : 
        MX2
      port map(A => \sample_in_buf[51]\, B => sample_4(2), S => 
        sample_val_delay, Y => \sample_in_buf_989[69]\);
    
    \loop_all_sample.14.loop_all_chanel.6.sample_in_buf[21]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_205[21]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[21]\);
    
    \loop_all_sample.9.loop_all_chanel.5.sample_in_buf[44]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_533[44]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[44]\);
    
    \loop_all_sample.11.loop_all_chanel.5.sample_in_buf[42]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_405[42]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[42]\);
    
    \loop_all_sample.9.loop_all_chanel.2.sample_in_buf_RNO[98]\ : 
        MX2
      port map(A => \sample_in_buf[80]\, B => sample_2(9), S => 
        sample_val_delay, Y => \sample_in_buf_557[98]\);
    
    \loop_all_sample.10.loop_all_chanel.4.sample_in_buf_RNO[61]\ : 
        MX2
      port map(A => \sample_in_buf[43]\, B => sample_4(10), S => 
        sample_val_delay, Y => \sample_in_buf_477[61]\);
    
    \chanel_more.all_chanel.1.all_bit.8.sample_out_s2[135]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[117]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_133);
    
    \loop_all_sample.9.loop_all_chanel.6.sample_in_buf[26]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_525[26]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[26]\);
    
    \chanel_more.all_chanel.1.all_bit.9.sample_out_s2[134]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[116]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_132);
    
    \loop_all_sample.11.loop_all_chanel.7.sample_in_buf_RNO[6]\ : 
        MX2
      port map(A => \sample_in_buf[132]\, B => sample_7(11), S
         => sample_val_delay, Y => \sample_in_buf_389[6]\);
    
    \loop_all_sample.1.loop_all_chanel.6.sample_in_buf_RNO[34]\ : 
        MX2
      port map(A => \sample_in_buf[16]\, B => sample_6(1), S => 
        sample_val_delay, Y => \sample_in_buf_1037[34]\);
    
    \loop_all_sample.3.loop_all_chanel.3.sample_in_buf[86]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_933[86]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[86]\);
    
    \chanel_more.all_chanel.6.all_bit.1.sample_out_s2[52]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[34]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[52]\);
    
    \chanel_HIGH.6.sample_out_s2[11]\ : DFN1E1C0
      port map(D => \sample_out_s[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[11]\);
    
    \loop_all_sample.11.loop_all_chanel.2.sample_in_buf_RNO[96]\ : 
        MX2
      port map(A => \sample_in_buf[78]\, B => sample_2(11), S => 
        sample_val_delay, Y => \sample_in_buf_429[96]\);
    
    \chanel_more.all_chanel.1.all_bit.5.sample_out_s2[138]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[120]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_136);
    
    \loop_all_sample.2.loop_all_chanel.7.sample_in_buf_RNO[15]\ : 
        MX2
      port map(A => \sample_in_buf[141]\, B => sample_7(2), S => 
        sample_val_delay, Y => \sample_in_buf_965[15]\);
    
    \loop_all_sample.13.loop_all_chanel.2.sample_in_buf[94]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_301[94]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[94]\);
    
    \loop_all_sample.17.loop_all_chanel.1.sample_in_buf[108]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_53[108]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[108]\);
    
    \loop_all_sample.0.loop_all_chanel.6.sample_in_buf_RNO[35]\ : 
        MX2
      port map(A => \sample_in_buf[17]\, B => sample_6(0), S => 
        sample_val_delay, Y => \sample_in_buf_1101[35]\);
    
    \loop_all_sample.4.loop_all_chanel.0.sample_in_buf_RNO[139]\ : 
        MX2
      port map(A => \sample_in_buf[121]\, B => sample_0(4), S => 
        sample_val_delay, Y => \sample_in_buf_893[139]\);
    
    \loop_all_sample.0.loop_all_chanel.3.sample_in_buf[89]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1125[89]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[89]\);
    
    \chanel_more.all_chanel.5.all_bit.9.sample_out_s2[62]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[44]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[62]\);
    
    \loop_all_sample.11.loop_all_chanel.2.sample_in_buf[96]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_429[96]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[96]\);
    
    \loop_all_sample.1.loop_all_chanel.3.sample_in_buf[88]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1061[88]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[88]\);
    
    \chanel_more.all_chanel.4.all_bit.11.sample_out_s2[78]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[60]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[78]\);
    
    \chanel_HIGH.15.sample_out_s2[2]\ : DFN1E1C0
      port map(D => \sample_out_s[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[2]\);
    
    \loop_all_sample.0.loop_all_chanel.5.sample_in_buf_RNO[53]\ : 
        MX2
      port map(A => \sample_in_buf[35]\, B => sample_5(0), S => 
        sample_val_delay, Y => \sample_in_buf_1109[53]\);
    
    \loop_all_sample.6.loop_all_chanel.4.sample_in_buf[65]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_733[65]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[65]\);
    
    \loop_all_sample.7.loop_all_chanel.7.sample_in_buf_RNO[10]\ : 
        MX2
      port map(A => \sample_in_buf[136]\, B => sample_7(7), S => 
        sample_val_delay, Y => \sample_in_buf_645[10]\);
    
    \loop_all_sample.17.loop_all_chanel.4.sample_in_buf[54]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_29[54]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[54]\);
    
    \loop_all_sample.4.loop_all_chanel.1.sample_in_buf_RNO[121]\ : 
        MX2
      port map(A => \sample_in_buf[103]\, B => sample_1(4), S => 
        sample_val_delay, Y => \sample_in_buf_885[121]\);
    
    \loop_all_sample.13.loop_all_chanel.6.sample_in_buf[22]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_269[22]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[22]\);
    
    \loop_all_sample.17.loop_all_chanel.2.sample_in_buf_RNO[90]\ : 
        MX2
      port map(A => \sample_in_buf[72]\, B => sample_2(15), S => 
        sample_val_delay, Y => \sample_in_buf_45[90]\);
    
    \loop_all_sample.11.loop_all_chanel.6.sample_in_buf_RNO[24]\ : 
        MX2
      port map(A => \sample_in_buf[6]\, B => sample_6(11), S => 
        sample_val_delay, Y => \sample_in_buf_397[24]\);
    
    \loop_all_sample.1.loop_all_chanel.7.sample_in_buf_RNO[16]\ : 
        MX2
      port map(A => \sample_in_buf[142]\, B => sample_7(1), S => 
        sample_val_delay, Y => \sample_in_buf_1029[16]\);
    
    \loop_all_sample.6.loop_all_chanel.7.sample_in_buf[11]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_709[11]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[11]\);
    
    \chanel_more.all_chanel.6.all_bit.8.sample_out_s2[45]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[27]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[45]\);
    
    \loop_all_sample.7.loop_all_chanel.0.sample_in_buf_RNO[136]\ : 
        MX2
      port map(A => \sample_in_buf[118]\, B => sample_0(7), S => 
        sample_val_delay, Y => \sample_in_buf_701[136]\);
    
    \chanel_more.all_chanel.3.all_bit.10.sample_out_s2[97]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[79]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[97]\);
    
    \loop_all_sample.4.loop_all_chanel.5.sample_in_buf_RNO[49]\ : 
        MX2
      port map(A => \sample_in_buf[31]\, B => sample_5(4), S => 
        sample_val_delay, Y => \sample_in_buf_853[49]\);
    
    \chanel_more.all_chanel.1.all_bit.13.sample_out_s2[130]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[112]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_128);
    
    \loop_all_sample.13.loop_all_chanel.5.sample_in_buf_RNO[40]\ : 
        MX2
      port map(A => \sample_in_buf[22]\, B => sample_5(13), S => 
        sample_val_delay, Y => \sample_in_buf_277[40]\);
    
    \loop_all_sample.17.loop_all_chanel.3.sample_in_buf[72]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_37[72]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[72]\);
    
    \chanel_more.all_chanel.6.all_bit.12.sample_out_s2[41]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[23]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[41]\);
    
    \chanel_more.all_chanel.4.all_bit.4.sample_out_s2[85]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[67]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[85]\);
    
    \loop_all_sample.5.loop_all_chanel.1.sample_in_buf[120]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_821[120]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[120]\);
    
    \loop_all_sample.11.loop_all_chanel.4.sample_in_buf_RNO[60]\ : 
        MX2
      port map(A => \sample_in_buf[42]\, B => sample_4(11), S => 
        sample_val_delay, Y => \sample_in_buf_413[60]\);
    
    \loop_all_sample.0.loop_all_chanel.1.sample_in_buf_RNO[125]\ : 
        MX2
      port map(A => \sample_in_buf[107]\, B => sample_1(0), S => 
        sample_val_delay, Y => \sample_in_buf_1141[125]\);
    
    \loop_all_sample.7.loop_all_chanel.2.sample_in_buf[100]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_685[100]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[100]\);
    
    \loop_all_sample.9.loop_all_chanel.7.sample_in_buf[8]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_517[8]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[8]\);
    
    \chanel_more.all_chanel.2.all_bit.7.sample_out_s2[118]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[100]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[118]\);
    
    \chanel_HIGH.9.sample_out_s2[8]\ : DFN1E1C0
      port map(D => \sample_out_s[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[8]\);
    
    \loop_all_sample.6.loop_all_chanel.5.sample_in_buf[47]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_725[47]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[47]\);
    
    \loop_all_sample.13.loop_all_chanel.4.sample_in_buf[58]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_285[58]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[58]\);
    
    \chanel_more.all_chanel.4.all_bit.5.sample_out_s2[84]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[66]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[84]\);
    
    \loop_all_sample.4.loop_all_chanel.2.sample_in_buf[103]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_877[103]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[103]\);
    
    \loop_all_sample.1.loop_all_chanel.7.sample_in_buf[16]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1029[16]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[16]\);
    
    \chanel_HIGH.7.sample_out_s2[10]\ : DFN1E1C0
      port map(D => \sample_out_s[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[10]\);
    
    \loop_all_sample.13.loop_all_chanel.7.sample_in_buf_RNO[4]\ : 
        MX2
      port map(A => \sample_in_buf[130]\, B => sample_7(13), S
         => sample_val_delay, Y => \sample_in_buf_261[4]\);
    
    \loop_all_sample.11.loop_all_chanel.7.sample_in_buf[6]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_389[6]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[6]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \loop_all_sample.1.loop_all_chanel.3.sample_in_buf_RNO[88]\ : 
        MX2
      port map(A => \sample_in_buf[70]\, B => sample_3(1), S => 
        sample_val_delay, Y => \sample_in_buf_1061[88]\);
    
    \loop_all_sample.13.loop_all_chanel.4.sample_in_buf_RNO[58]\ : 
        MX2
      port map(A => \sample_in_buf[40]\, B => sample_4(13), S => 
        sample_val_delay, Y => \sample_in_buf_285[58]\);
    
    \chanel_more.all_chanel.1.all_bit.4.sample_out_s2[139]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[121]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_137);
    
    \chanel_more.all_chanel.7.all_bit.6.sample_out_s2[29]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[11]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[29]\);
    
    \loop_all_sample.2.loop_all_chanel.2.sample_in_buf_RNO[105]\ : 
        MX2
      port map(A => \sample_in_buf[87]\, B => sample_2(2), S => 
        sample_val_delay, Y => \sample_in_buf_1005[105]\);
    
    \loop_all_sample.10.loop_all_chanel.2.sample_in_buf[97]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_493[97]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[97]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \loop_all_sample.2.loop_all_chanel.5.sample_in_buf_RNO[51]\ : 
        MX2
      port map(A => \sample_in_buf[33]\, B => sample_5(2), S => 
        sample_val_delay, Y => \sample_in_buf_981[51]\);
    
    \loop_all_sample.17.loop_all_chanel.5.sample_in_buf[36]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_21[36]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[36]\);
    
    \loop_all_sample.17.loop_all_chanel.3.sample_in_buf_RNO[72]\ : 
        MX2
      port map(A => \sample_in_buf[54]\, B => sample_3(15), S => 
        sample_val_delay, Y => \sample_in_buf_37[72]\);
    
    \chanel_more.all_chanel.2.all_bit.9.sample_out_s2[116]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[98]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[116]\);
    
    \loop_all_sample.7.loop_all_chanel.1.sample_in_buf_RNO[118]\ : 
        MX2
      port map(A => \sample_in_buf[100]\, B => sample_1(7), S => 
        sample_val_delay, Y => \sample_in_buf_693[118]\);
    
    \chanel_more.all_chanel.2.all_bit.10.sample_out_s2[115]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[97]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[115]\);
    
    \chanel_more.all_chanel.3.all_bit.6.sample_out_s2[101]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[83]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[101]\);
    
    \loop_all_sample.9.loop_all_chanel.4.sample_in_buf[62]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_541[62]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[62]\);
    
    \loop_all_sample.14.loop_all_chanel.0.sample_in_buf[129]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_253[129]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[129]\);
    
    \loop_all_sample.7.loop_all_chanel.0.sample_in_buf[136]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_701[136]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[136]\);
    
    \chanel_more.all_chanel.4.all_bit.0.sample_out_s2[89]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[71]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[89]\);
    
    \loop_all_sample.3.loop_all_chanel.2.sample_in_buf[104]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_941[104]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[104]\);
    
    \loop_all_sample.5.loop_all_chanel.2.sample_in_buf_RNO[102]\ : 
        MX2
      port map(A => \sample_in_buf[84]\, B => sample_2(5), S => 
        sample_val_delay, Y => \sample_in_buf_813[102]\);
    
    \loop_all_sample.4.loop_all_chanel.1.sample_in_buf[121]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_885[121]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[121]\);
    
    \chanel_more.all_chanel.6.all_bit.11.sample_out_s2[42]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[24]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[42]\);
    
    \loop_all_sample.10.loop_all_chanel.5.sample_in_buf[43]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_469[43]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[43]\);
    
    \chanel_more.all_chanel.5.all_bit.0.sample_out_s2[71]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[53]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[71]\);
    
    \loop_all_sample.11.loop_all_chanel.0.sample_in_buf_RNO[132]\ : 
        MX2
      port map(A => \sample_in_buf[114]\, B => sample_0(11), S
         => sample_val_delay, Y => \sample_in_buf_445[132]\);
    
    \chanel_more.all_chanel.6.all_bit.6.sample_out_s2[47]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[29]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[47]\);
    
    \loop_all_sample.12.loop_all_chanel.2.sample_in_buf[95]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_365[95]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[95]\);
    
    \chanel_more.all_chanel.7.all_bit.1.sample_out_s2[34]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[16]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[34]\);
    
    \loop_all_sample.6.loop_all_chanel.2.sample_in_buf[101]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_749[101]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[101]\);
    
    \loop_all_sample.9.loop_all_chanel.1.sample_in_buf_RNO[116]\ : 
        MX2
      port map(A => \sample_in_buf[98]\, B => sample_1(9), S => 
        sample_val_delay, Y => \sample_in_buf_565[116]\);
    
    \loop_all_sample.4.loop_all_chanel.2.sample_in_buf_RNO[103]\ : 
        MX2
      port map(A => \sample_in_buf[85]\, B => sample_2(4), S => 
        sample_val_delay, Y => \sample_in_buf_877[103]\);
    
    \loop_all_sample.10.loop_all_chanel.1.sample_in_buf_RNO[115]\ : 
        MX2
      port map(A => \sample_in_buf[97]\, B => sample_1(10), S => 
        sample_val_delay, Y => \sample_in_buf_501[115]\);
    
    \loop_all_sample.5.loop_all_chanel.5.sample_in_buf_RNO[48]\ : 
        MX2
      port map(A => \sample_in_buf[30]\, B => sample_5(5), S => 
        sample_val_delay, Y => \sample_in_buf_789[48]\);
    
    \loop_all_sample.3.loop_all_chanel.2.sample_in_buf_RNO[104]\ : 
        MX2
      port map(A => \sample_in_buf[86]\, B => sample_2(3), S => 
        sample_val_delay, Y => \sample_in_buf_941[104]\);
    
    \chanel_more.all_chanel.7.all_bit.15.sample_out_s2[20]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[20]\);
    
    \loop_all_sample.2.loop_all_chanel.1.sample_in_buf[123]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1013[123]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[123]\);
    
    \chanel_HIGH.13.sample_out_s2[4]\ : DFN1E1C0
      port map(D => \sample_out_s[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[4]\);
    
    \loop_all_sample.10.loop_all_chanel.6.sample_in_buf[25]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_461[25]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[25]\);
    
    \chanel_more.all_chanel.3.all_bit.13.sample_out_s2[94]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[76]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[94]\);
    
    \loop_all_sample.3.loop_all_chanel.1.sample_in_buf_RNO[122]\ : 
        MX2
      port map(A => \sample_in_buf[104]\, B => sample_1(3), S => 
        sample_val_delay, Y => \sample_in_buf_949[122]\);
    
    \loop_all_sample.2.loop_all_chanel.1.sample_in_buf_RNO[123]\ : 
        MX2
      port map(A => \sample_in_buf[105]\, B => sample_1(2), S => 
        sample_val_delay, Y => \sample_in_buf_1013[123]\);
    
    \loop_all_sample.3.loop_all_chanel.0.sample_in_buf_RNO[140]\ : 
        MX2
      port map(A => \sample_in_buf[122]\, B => sample_0(3), S => 
        sample_val_delay, Y => \sample_in_buf_957[140]\);
    
    \loop_all_sample.7.loop_all_chanel.6.sample_in_buf_RNO[28]\ : 
        MX2
      port map(A => \sample_in_buf[10]\, B => sample_6(7), S => 
        sample_val_delay, Y => \sample_in_buf_653[28]\);
    
    \loop_all_sample.8.loop_all_chanel.3.sample_in_buf_RNO[81]\ : 
        MX2
      port map(A => \sample_in_buf[63]\, B => sample_3(8), S => 
        sample_val_delay, Y => \sample_in_buf_613[81]\);
    
    \loop_all_sample.14.loop_all_chanel.5.sample_in_buf_RNO[39]\ : 
        MX2
      port map(A => \sample_in_buf[21]\, B => sample_5(14), S => 
        sample_val_delay, Y => \sample_in_buf_213[39]\);
    
    \loop_all_sample.12.loop_all_chanel.7.sample_in_buf_RNO[5]\ : 
        MX2
      port map(A => \sample_in_buf[131]\, B => sample_7(12), S
         => sample_val_delay, Y => \sample_in_buf_325[5]\);
    
    \loop_all_sample.0.loop_all_chanel.2.sample_in_buf_RNO[107]\ : 
        MX2
      port map(A => \sample_in_buf[89]\, B => sample_2(0), S => 
        sample_val_delay, Y => \sample_in_buf_1133[107]\);
    
    \chanel_more.all_chanel.1.all_bit.15.sample_out_s2[128]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[110]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_126);
    
    \loop_all_sample.8.loop_all_chanel.1.sample_in_buf[117]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_629[117]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[117]\);
    
    \loop_all_sample.11.loop_all_chanel.1.sample_in_buf_RNO[114]\ : 
        MX2
      port map(A => \sample_in_buf[96]\, B => sample_1(11), S => 
        sample_val_delay, Y => \sample_in_buf_437[114]\);
    
    \loop_all_sample.5.loop_all_chanel.3.sample_in_buf_RNO[84]\ : 
        MX2
      port map(A => \sample_in_buf[66]\, B => sample_3(5), S => 
        sample_val_delay, Y => \sample_in_buf_805[84]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \chanel_more.all_chanel.6.all_bit.3.sample_out_s2[50]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[32]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[50]\);
    
    \loop_all_sample.2.loop_all_chanel.5.sample_in_buf[51]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_981[51]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[51]\);
    
    \chanel_more.all_chanel.7.all_bit.7.sample_out_s2[28]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[10]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[28]\);
    
    \chanel_more.all_chanel.2.all_bit.15.sample_out_s2[110]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[92]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[110]\);
    
    \loop_all_sample.8.loop_all_chanel.5.sample_in_buf[45]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_597[45]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[45]\);
    
    \loop_all_sample.9.loop_all_chanel.7.sample_in_buf_RNO[8]\ : 
        MX2
      port map(A => \sample_in_buf[134]\, B => sample_7(9), S => 
        sample_val_delay, Y => \sample_in_buf_517[8]\);
    
    \loop_all_sample.4.loop_all_chanel.6.sample_in_buf_RNO[31]\ : 
        MX2
      port map(A => \sample_in_buf[13]\, B => sample_6(4), S => 
        sample_val_delay, Y => \sample_in_buf_845[31]\);
    
    \loop_all_sample.8.loop_all_chanel.5.sample_in_buf_RNO[45]\ : 
        MX2
      port map(A => \sample_in_buf[27]\, B => sample_5(8), S => 
        sample_val_delay, Y => \sample_in_buf_597[45]\);
    
    \loop_all_sample.11.loop_all_chanel.1.sample_in_buf[114]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_437[114]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[114]\);
    
    \loop_all_sample.2.loop_all_chanel.0.sample_in_buf[141]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1021[141]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[141]\);
    
    \loop_all_sample.14.loop_all_chanel.4.sample_in_buf[57]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_221[57]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[57]\);
    
    IIR_CEL_CTRLR_v2_DATAFLOW_1 : IIR_CEL_CTRLR_v2_DATAFLOW
      port map(alu_ctrl(2) => \alu_ctrl[2]\, alu_ctrl(1) => 
        \alu_ctrl[1]\, alu_ctrl(0) => \alu_ctrl[0]\, S(8) => 
        \S[8]\, S_i_0(33) => \S_i_0[33]\, alu_sel_coeff(4) => 
        \alu_sel_coeff[4]\, alu_sel_coeff(3) => 
        \alu_sel_coeff[3]\, alu_sel_coeff(2) => 
        \alu_sel_coeff[2]\, alu_sel_coeff(1) => 
        \alu_sel_coeff[1]\, alu_sel_coeff(0) => 
        \alu_sel_coeff[0]\, alu_sel_coeff_0_2 => 
        \alu_sel_coeff_0[2]\, alu_sel_coeff_0_0 => 
        \alu_sel_coeff_0[0]\, waddr_previous(1) => 
        \waddr_previous[1]\, waddr_previous(0) => 
        \waddr_previous[0]\, sample_0(14) => sample_0(14), 
        sample_0(13) => sample_0(13), sample_0(12) => 
        sample_0(12), sample_0(11) => sample_0(11), sample_0(10)
         => sample_0(10), sample_0(9) => sample_0(9), sample_0(8)
         => sample_0(8), sample_0(7) => sample_0(7), sample_0(6)
         => sample_0(6), sample_0(5) => sample_0(5), sample_0(4)
         => sample_0(4), sample_0(3) => sample_0(3), sample_0(2)
         => sample_0(2), sample_0(1) => sample_0(1), sample_0(0)
         => sample_0(0), sample_in_buf(143) => 
        \sample_in_buf[143]\, sample_in_buf(142) => 
        \sample_in_buf[142]\, sample_in_buf(141) => 
        \sample_in_buf[141]\, sample_in_buf(140) => 
        \sample_in_buf[140]\, sample_in_buf(139) => 
        \sample_in_buf[139]\, sample_in_buf(138) => 
        \sample_in_buf[138]\, sample_in_buf(137) => 
        \sample_in_buf[137]\, sample_in_buf(136) => 
        \sample_in_buf[136]\, sample_in_buf(135) => 
        \sample_in_buf[135]\, sample_in_buf(134) => 
        \sample_in_buf[134]\, sample_in_buf(133) => 
        \sample_in_buf[133]\, sample_in_buf(132) => 
        \sample_in_buf[132]\, sample_in_buf(131) => 
        \sample_in_buf[131]\, sample_in_buf(130) => 
        \sample_in_buf[130]\, sample_in_buf(129) => 
        \sample_in_buf[129]\, ram_sel_Wdata(1) => 
        \ram_sel_Wdata[1]\, ram_sel_Wdata(0) => 
        \ram_sel_Wdata[0]\, sample_out_s_0 => \sample_out_s[0]\, 
        sample_out_s_1 => \sample_out_s[1]\, sample_out_s_3 => 
        \sample_out_s[3]\, sample_out_s_2 => \sample_out_s[2]\, 
        sample_out_s_10 => \sample_out_s[10]\, sample_out_s_15
         => \sample_out_s[15]\, sample_out_s_14 => 
        \sample_out_s[14]\, sample_out_s_13 => \sample_out_s[13]\, 
        sample_out_s_12 => \sample_out_s[12]\, sample_out_s_11
         => \sample_out_s[11]\, sample_out_s_9 => 
        \sample_out_s[9]\, sample_out_s_8 => \sample_out_s[8]\, 
        sample_out_s_7 => \sample_out_s[7]\, sample_out_s_6 => 
        \sample_out_s[6]\, sample_out_s_5 => \sample_out_s[5]\, 
        sample_out_s_4 => \sample_out_s[4]\, sample_in_s_1(17)
         => \sample_in_s_1[17]\, in_sel_src(1) => \in_sel_src[1]\, 
        in_sel_src(0) => \in_sel_src[0]\, raddr_rst => raddr_rst, 
        raddr_add1 => raddr_add1, ram_write => ram_write, 
        IIR_CEL_CTRLR_v2_DATAFLOW_GND => IIR_CEL_CTRLR_v2_GND, 
        IIR_CEL_CTRLR_v2_DATAFLOW_VCC => IIR_CEL_CTRLR_v2_VCC, 
        ram_write_i => ram_write_i, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, sample_val_delay => sample_val_delay, 
        alu_sel_input => alu_sel_input);
    
    sample_out_val : DFN1C0
      port map(D => \sample_out_val_s2\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_filter_v2_out_val);
    
    \loop_all_sample.8.loop_all_chanel.3.sample_in_buf[81]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_613[81]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[81]\);
    
    \loop_all_sample.17.loop_all_chanel.4.sample_in_buf_RNO[54]\ : 
        MX2
      port map(A => \sample_in_buf[36]\, B => sample_4(15), S => 
        sample_val_delay, Y => \sample_in_buf_29[54]\);
    
    \loop_all_sample.4.loop_all_chanel.3.sample_in_buf[85]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_869[85]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[85]\);
    
    \loop_all_sample.3.loop_all_chanel.4.sample_in_buf[68]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_925[68]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[68]\);
    
    \loop_all_sample.10.loop_all_chanel.7.sample_in_buf_RNO[7]\ : 
        MX2
      port map(A => \sample_in_buf[133]\, B => sample_7(10), S
         => sample_val_delay, Y => \sample_in_buf_453[7]\);
    
    \loop_all_sample.10.loop_all_chanel.4.sample_in_buf[61]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_477[61]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[61]\);
    
    \loop_all_sample.10.loop_all_chanel.3.sample_in_buf[79]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_485[79]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[79]\);
    
    \chanel_more.all_chanel.4.all_bit.15.sample_out_s2[74]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[56]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[74]\);
    
    \chanel_more.all_chanel.2.all_bit.5.sample_out_s2[120]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[102]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[120]\);
    
    \chanel_more.all_chanel.2.all_bit.14.sample_out_s2[111]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[93]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[111]\);
    
    \chanel_more.all_chanel.2.all_bit.6.sample_out_s2[119]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[101]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[119]\);
    
    \loop_all_sample.11.loop_all_chanel.0.sample_in_buf[132]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_445[132]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[132]\);
    
    \chanel_more.all_chanel.7.all_bit.13.sample_out_s2[22]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[22]\);
    
    \loop_all_sample.6.loop_all_chanel.5.sample_in_buf_RNO[47]\ : 
        MX2
      port map(A => \sample_in_buf[29]\, B => sample_5(6), S => 
        sample_val_delay, Y => \sample_in_buf_725[47]\);
    
    \loop_all_sample.17.loop_all_chanel.0.sample_in_buf_RNO[126]\ : 
        MX2
      port map(A => \sample_in_buf[108]\, B => sample_0(15), S
         => sample_val_delay, Y => \sample_in_buf_61[126]\);
    
    \loop_all_sample.6.loop_all_chanel.6.sample_in_buf[29]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_717[29]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[29]\);
    
    \loop_all_sample.1.loop_all_chanel.2.sample_in_buf_RNO[106]\ : 
        MX2
      port map(A => \sample_in_buf[88]\, B => sample_2(1), S => 
        sample_val_delay, Y => \sample_in_buf_1069[106]\);
    
    \loop_all_sample.0.loop_all_chanel.6.sample_in_buf[35]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1101[35]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[35]\);
    
    \chanel_more.all_chanel.3.all_bit.0.sample_out_s2[107]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[89]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[107]\);
    
    \loop_all_sample.4.loop_all_chanel.6.sample_in_buf[31]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_845[31]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[31]\);
    
    \chanel_more.all_chanel.4.all_bit.8.sample_out_s2[81]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[63]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[81]\);
    
    \chanel_more.all_chanel.6.all_bit.14.sample_out_s2[39]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[21]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[39]\);
    
    \loop_all_sample.12.loop_all_chanel.3.sample_in_buf_RNO[77]\ : 
        MX2
      port map(A => \sample_in_buf[59]\, B => sample_3(12), S => 
        sample_val_delay, Y => \sample_in_buf_357[77]\);
    
    \loop_all_sample.1.loop_all_chanel.5.sample_in_buf_RNO[52]\ : 
        MX2
      port map(A => \sample_in_buf[34]\, B => sample_5(1), S => 
        sample_val_delay, Y => \sample_in_buf_1045[52]\);
    
    \chanel_more.all_chanel.7.all_bit.14.sample_out_s2[21]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[21]\);
    
    \loop_all_sample.2.loop_all_chanel.2.sample_in_buf[105]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1005[105]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[105]\);
    
    \loop_all_sample.10.loop_all_chanel.6.sample_in_buf_RNO[25]\ : 
        MX2
      port map(A => \sample_in_buf[7]\, B => sample_6(10), S => 
        sample_val_delay, Y => \sample_in_buf_461[25]\);
    
    \chanel_more.all_chanel.3.all_bit.14.sample_out_s2[93]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[75]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[93]\);
    
    \loop_all_sample.2.loop_all_chanel.0.sample_in_buf_RNO[141]\ : 
        MX2
      port map(A => \sample_in_buf[123]\, B => sample_0(2), S => 
        sample_val_delay, Y => \sample_in_buf_1021[141]\);
    
    \loop_all_sample.3.loop_all_chanel.1.sample_in_buf[122]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_949[122]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[122]\);
    
    \chanel_more.all_chanel.4.all_bit.9.sample_out_s2[80]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[62]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[80]\);
    
    \chanel_more.all_chanel.4.all_bit.6.sample_out_s2[83]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[65]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[83]\);
    
    \loop_all_sample.13.loop_all_chanel.6.sample_in_buf_RNO[22]\ : 
        MX2
      port map(A => \sample_in_buf[4]\, B => sample_6(13), S => 
        sample_val_delay, Y => \sample_in_buf_269[22]\);
    
    \loop_all_sample.8.loop_all_chanel.6.sample_in_buf[27]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_589[27]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[27]\);
    
    \loop_all_sample.2.loop_all_chanel.3.sample_in_buf[87]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_997[87]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[87]\);
    
    \chanel_more.all_chanel.3.all_bit.15.sample_out_s2[92]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[74]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[92]\);
    
    \loop_all_sample.3.loop_all_chanel.3.sample_in_buf_RNO[86]\ : 
        MX2
      port map(A => \sample_in_buf[68]\, B => sample_3(3), S => 
        sample_val_delay, Y => \sample_in_buf_933[86]\);
    
    \chanel_more.all_chanel.6.all_bit.10.sample_out_s2[43]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[25]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[43]\);
    
    \loop_all_sample.6.loop_all_chanel.4.sample_in_buf_RNO[65]\ : 
        MX2
      port map(A => \sample_in_buf[47]\, B => sample_4(6), S => 
        sample_val_delay, Y => \sample_in_buf_733[65]\);
    
    \loop_all_sample.0.loop_all_chanel.0.sample_in_buf[143]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1149[143]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[143]\);
    
    \loop_all_sample.3.loop_all_chanel.0.sample_in_buf[140]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_957[140]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[140]\);
    
    \loop_all_sample.1.loop_all_chanel.4.sample_in_buf[70]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1053[70]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[70]\);
    
    \loop_all_sample.14.loop_all_chanel.2.sample_in_buf[93]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_237[93]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[93]\);
    
    \chanel_HIGH.14.sample_out_s2[3]\ : DFN1E1C0
      port map(D => \sample_out_s[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[3]\);
    
    \loop_all_sample.9.loop_all_chanel.1.sample_in_buf[116]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_565[116]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[116]\);
    
    \loop_all_sample.17.loop_all_chanel.2.sample_in_buf[90]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_45[90]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[90]\);
    
    \loop_all_sample.0.loop_all_chanel.2.sample_in_buf[107]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1133[107]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[107]\);
    
    \loop_all_sample.4.loop_all_chanel.4.sample_in_buf_RNO[67]\ : 
        MX2
      port map(A => \sample_in_buf[49]\, B => sample_4(4), S => 
        sample_val_delay, Y => \sample_in_buf_861[67]\);
    
    \loop_all_sample.8.loop_all_chanel.0.sample_in_buf[135]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_637[135]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[135]\);
    
    \chanel_more.all_chanel.5.all_bit.13.sample_out_s2[58]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[40]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[58]\);
    
    \chanel_HIGH.2.sample_out_s2[15]\ : DFN1E1C0
      port map(D => \sample_out_s[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[15]\);
    
    \chanel_more.all_chanel.4.all_bit.10.sample_out_s2[79]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[61]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[79]\);
    
    \loop_all_sample.12.loop_all_chanel.2.sample_in_buf_RNO[95]\ : 
        MX2
      port map(A => \sample_in_buf[77]\, B => sample_2(12), S => 
        sample_val_delay, Y => \sample_in_buf_365[95]\);
    
    \loop_all_sample.5.loop_all_chanel.5.sample_in_buf[48]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_789[48]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[48]\);
    
    \loop_all_sample.14.loop_all_chanel.7.sample_in_buf[3]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_197[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[3]\);
    
    \chanel_more.all_chanel.7.all_bit.10.sample_out_s2[25]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[7]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[25]\);
    
    \loop_all_sample.12.loop_all_chanel.3.sample_in_buf[77]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_357[77]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[77]\);
    
    \chanel_more.all_chanel.3.all_bit.3.sample_out_s2[104]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[86]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[104]\);
    
    sample_out_val_s2 : DFN1C0
      port map(D => sample_out_val_s, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sample_out_val_s2\);
    
    \chanel_more.all_chanel.7.all_bit.9.sample_out_s2[26]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[8]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[26]\);
    
    \loop_all_sample.5.loop_all_chanel.6.sample_in_buf_RNO[30]\ : 
        MX2
      port map(A => \sample_in_buf[12]\, B => sample_6(5), S => 
        sample_val_delay, Y => \sample_in_buf_781[30]\);
    
    \loop_all_sample.14.loop_all_chanel.5.sample_in_buf[39]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_213[39]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[39]\);
    
    \chanel_more.all_chanel.2.all_bit.0.sample_out_s2[125]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[107]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[125]\);
    
    \chanel_more.all_chanel.2.all_bit.2.sample_out_s2[123]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[105]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[123]\);
    
    \chanel_more.all_chanel.3.all_bit.7.sample_out_s2[100]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[82]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[100]\);
    
    \loop_all_sample.4.loop_all_chanel.7.sample_in_buf_RNO[13]\ : 
        MX2
      port map(A => \sample_in_buf[139]\, B => sample_7(4), S => 
        sample_val_delay, Y => \sample_in_buf_837[13]\);
    
    \loop_all_sample.14.loop_all_chanel.6.sample_in_buf_RNO[21]\ : 
        MX2
      port map(A => \sample_in_buf[3]\, B => sample_6(14), S => 
        sample_val_delay, Y => \sample_in_buf_205[21]\);
    
    \chanel_more.all_chanel.2.all_bit.13.sample_out_s2[112]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[94]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[112]\);
    
    \loop_all_sample.9.loop_all_chanel.6.sample_in_buf_RNO[26]\ : 
        MX2
      port map(A => \sample_in_buf[8]\, B => sample_6(9), S => 
        sample_val_delay, Y => \sample_in_buf_525[26]\);
    
    \loop_all_sample.9.loop_all_chanel.3.sample_in_buf[80]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_549[80]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[80]\);
    
    \loop_all_sample.7.loop_all_chanel.7.sample_in_buf[10]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_645[10]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[10]\);
    
    \loop_all_sample.12.loop_all_chanel.1.sample_in_buf_RNO[113]\ : 
        MX2
      port map(A => \sample_in_buf[95]\, B => sample_1(12), S => 
        sample_val_delay, Y => \sample_in_buf_373[113]\);
    
    \chanel_HIGH.1.sample_out_s2[16]\ : DFN1E1C0
      port map(D => \sample_out_s[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[16]\);
    
    \loop_all_sample.8.loop_all_chanel.4.sample_in_buf_RNO[63]\ : 
        MX2
      port map(A => \sample_in_buf[45]\, B => sample_4(8), S => 
        sample_val_delay, Y => \sample_in_buf_605[63]\);
    
    \loop_all_sample.6.loop_all_chanel.7.sample_in_buf_RNO[11]\ : 
        MX2
      port map(A => \sample_in_buf[137]\, B => sample_7(6), S => 
        sample_val_delay, Y => \sample_in_buf_709[11]\);
    
    \loop_all_sample.14.loop_all_chanel.0.sample_in_buf_RNO[129]\ : 
        MX2
      port map(A => \sample_in_buf[111]\, B => sample_0(14), S
         => sample_val_delay, Y => \sample_in_buf_253[129]\);
    
    \chanel_HIGH.12.sample_out_s2[5]\ : DFN1E1C0
      port map(D => \sample_out_s[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[5]\);
    
    \loop_all_sample.3.loop_all_chanel.6.sample_in_buf[32]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_909[32]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[32]\);
    
    \loop_all_sample.17.loop_all_chanel.5.sample_in_buf_RNO[36]\ : 
        MX2
      port map(A => \sample_in_buf[18]\, B => sample_5(15), S => 
        sample_val_delay, Y => \sample_in_buf_21[36]\);
    
    \chanel_more.all_chanel.5.all_bit.8.sample_out_s2[63]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[45]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[63]\);
    
    \loop_all_sample.8.loop_all_chanel.7.sample_in_buf_RNO[9]\ : 
        MX2
      port map(A => \sample_in_buf[135]\, B => sample_7(8), S => 
        sample_val_delay, Y => \sample_in_buf_581[9]\);
    
    \loop_all_sample.5.loop_all_chanel.7.sample_in_buf_RNO[12]\ : 
        MX2
      port map(A => \sample_in_buf[138]\, B => sample_7(5), S => 
        sample_val_delay, Y => \sample_in_buf_773[12]\);
    
    \loop_all_sample.1.loop_all_chanel.4.sample_in_buf_RNO[70]\ : 
        MX2
      port map(A => \sample_in_buf[52]\, B => sample_4(1), S => 
        sample_val_delay, Y => \sample_in_buf_1053[70]\);
    
    \loop_all_sample.7.loop_all_chanel.6.sample_in_buf[28]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_653[28]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[28]\);
    
    \loop_all_sample.13.loop_all_chanel.3.sample_in_buf[76]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_293[76]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[76]\);
    
    \loop_all_sample.17.loop_all_chanel.6.sample_in_buf[18]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_13[18]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[18]\);
    
    \loop_all_sample.0.loop_all_chanel.3.sample_in_buf_RNO[89]\ : 
        MX2
      port map(A => \sample_in_buf[71]\, B => sample_3(0), S => 
        sample_val_delay, Y => \sample_in_buf_1125[89]\);
    
    \chanel_more.all_chanel.2.all_bit.11.sample_out_s2[114]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[96]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[114]\);
    
    \loop_all_sample.12.loop_all_chanel.1.sample_in_buf[113]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_373[113]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[113]\);
    
    \loop_all_sample.0.loop_all_chanel.4.sample_in_buf_RNO[71]\ : 
        MX2
      port map(A => \sample_in_buf[53]\, B => sample_4(0), S => 
        sample_val_delay, Y => \sample_in_buf_1117[71]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \loop_all_sample.13.loop_all_chanel.1.sample_in_buf[112]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_309[112]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[112]\);
    
    \chanel_more.all_chanel.6.all_bit.9.sample_out_s2[44]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[26]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[44]\);
    
    \chanel_more.all_chanel.2.all_bit.1.sample_out_s2[124]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[106]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[124]\);
    
    \loop_all_sample.12.loop_all_chanel.4.sample_in_buf[59]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_349[59]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[59]\);
    
    \loop_all_sample.8.loop_all_chanel.7.sample_in_buf[9]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_581[9]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[9]\);
    
    \chanel_HIGH.5.sample_out_s2[12]\ : DFN1E1C0
      port map(D => \sample_out_s[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[12]\);
    
    \loop_all_sample.5.loop_all_chanel.0.sample_in_buf[138]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_829[138]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[138]\);
    
    
        \loop_all_sample.17.loop_all_chanel.0.sample_in_buf_RNIF75G[126]\ : 
        MX2
      port map(A => \sample_in_buf[128]\, B => sample_0(15), S
         => sample_val_delay, Y => \sample_in_s_1[17]\);
    
    \loop_all_sample.3.loop_all_chanel.5.sample_in_buf[50]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_917[50]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[50]\);
    
    \loop_all_sample.0.loop_all_chanel.1.sample_in_buf[125]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1141[125]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[125]\);
    
    \loop_all_sample.9.loop_all_chanel.2.sample_in_buf[98]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_557[98]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[98]\);
    
    \loop_all_sample.6.loop_all_chanel.0.sample_in_buf[137]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_765[137]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[137]\);
    
    \loop_all_sample.3.loop_all_chanel.5.sample_in_buf_RNO[50]\ : 
        MX2
      port map(A => \sample_in_buf[32]\, B => sample_5(3), S => 
        sample_val_delay, Y => \sample_in_buf_917[50]\);
    
    \loop_all_sample.1.loop_all_chanel.1.sample_in_buf[124]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1077[124]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[124]\);
    
    \loop_all_sample.14.loop_all_chanel.3.sample_in_buf_RNO[75]\ : 
        MX2
      port map(A => \sample_in_buf[57]\, B => sample_3(14), S => 
        sample_val_delay, Y => \sample_in_buf_229[75]\);
    
    \chanel_HIGH.4.sample_out_s2[13]\ : DFN1E1C0
      port map(D => \sample_out_s[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[13]\);
    
    \chanel_HIGH.0.sample_out_s2[17]\ : DFN1E1C0
      port map(D => \sample_out_s[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[17]\);
    
    \loop_all_sample.7.loop_all_chanel.4.sample_in_buf[64]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_669[64]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[64]\);
    
    \chanel_more.all_chanel.1.all_bit.1.sample_out_s2[142]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[124]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_140);
    
    \loop_all_sample.6.loop_all_chanel.6.sample_in_buf_RNO[29]\ : 
        MX2
      port map(A => \sample_in_buf[11]\, B => sample_6(6), S => 
        sample_val_delay, Y => \sample_in_buf_717[29]\);
    
    \loop_all_sample.14.loop_all_chanel.4.sample_in_buf_RNO[57]\ : 
        MX2
      port map(A => \sample_in_buf[39]\, B => sample_4(14), S => 
        sample_val_delay, Y => \sample_in_buf_221[57]\);
    
    \loop_all_sample.12.loop_all_chanel.6.sample_in_buf_RNO[23]\ : 
        MX2
      port map(A => \sample_in_buf[5]\, B => sample_6(12), S => 
        sample_val_delay, Y => \sample_in_buf_333[23]\);
    
    \chanel_more.all_chanel.5.all_bit.4.sample_out_s2[67]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[49]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[67]\);
    
    \chanel_more.all_chanel.3.all_bit.9.sample_out_s2[98]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[80]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[98]\);
    
    \loop_all_sample.7.loop_all_chanel.5.sample_in_buf[46]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_661[46]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[46]\);
    
    \loop_all_sample.9.loop_all_chanel.0.sample_in_buf[134]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_573[134]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[134]\);
    
    \chanel_more.all_chanel.4.all_bit.3.sample_out_s2[86]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[68]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[86]\);
    
    \loop_all_sample.5.loop_all_chanel.7.sample_in_buf[12]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_773[12]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[12]\);
    
    \loop_all_sample.4.loop_all_chanel.7.sample_in_buf[13]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_837[13]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[13]\);
    
    \loop_all_sample.2.loop_all_chanel.4.sample_in_buf[69]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_989[69]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[69]\);
    
    \loop_all_sample.12.loop_all_chanel.0.sample_in_buf[131]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_381[131]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[131]\);
    
    \loop_all_sample.4.loop_all_chanel.5.sample_in_buf[49]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_853[49]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[49]\);
    
    \loop_all_sample.11.loop_all_chanel.6.sample_in_buf[24]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_397[24]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[24]\);
    
    \loop_all_sample.3.loop_all_chanel.7.sample_in_buf_RNO[14]\ : 
        MX2
      port map(A => \sample_in_buf[140]\, B => sample_7(3), S => 
        sample_val_delay, Y => \sample_in_buf_901[14]\);
    
    \loop_all_sample.1.loop_all_chanel.0.sample_in_buf[142]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1085[142]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[142]\);
    
    \loop_all_sample.8.loop_all_chanel.4.sample_in_buf[63]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_605[63]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[63]\);
    
    \loop_all_sample.10.loop_all_chanel.1.sample_in_buf[115]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_501[115]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[115]\);
    
    \loop_all_sample.0.loop_all_chanel.4.sample_in_buf[71]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1117[71]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[71]\);
    
    \loop_all_sample.4.loop_all_chanel.3.sample_in_buf_RNO[85]\ : 
        MX2
      port map(A => \sample_in_buf[67]\, B => sample_3(4), S => 
        sample_val_delay, Y => \sample_in_buf_869[85]\);
    
    \loop_all_sample.13.loop_all_chanel.3.sample_in_buf_RNO[76]\ : 
        MX2
      port map(A => \sample_in_buf[58]\, B => sample_3(13), S => 
        sample_val_delay, Y => \sample_in_buf_293[76]\);
    
    \loop_all_sample.14.loop_all_chanel.1.sample_in_buf[111]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_245[111]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[111]\);
    
    \chanel_more.all_chanel.3.all_bit.5.sample_out_s2[102]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[84]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[102]\);
    
    \loop_all_sample.2.loop_all_chanel.7.sample_in_buf[15]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_965[15]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[15]\);
    
    \loop_all_sample.14.loop_all_chanel.7.sample_in_buf_RNO[3]\ : 
        MX2
      port map(A => \sample_in_buf[129]\, B => sample_7(14), S
         => sample_val_delay, Y => \sample_in_buf_197[3]\);
    
    \chanel_more.all_chanel.7.all_bit.4.sample_out_s2[31]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[13]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[31]\);
    
    \loop_all_sample.7.loop_all_chanel.2.sample_in_buf_RNO[100]\ : 
        MX2
      port map(A => \sample_in_buf[82]\, B => sample_2(7), S => 
        sample_val_delay, Y => \sample_in_buf_685[100]\);
    
    \loop_all_sample.8.loop_all_chanel.0.sample_in_buf_RNO[135]\ : 
        MX2
      port map(A => \sample_in_buf[117]\, B => sample_0(8), S => 
        sample_val_delay, Y => \sample_in_buf_637[135]\);
    
    \loop_all_sample.7.loop_all_chanel.5.sample_in_buf_RNO[46]\ : 
        MX2
      port map(A => \sample_in_buf[28]\, B => sample_5(7), S => 
        sample_val_delay, Y => \sample_in_buf_661[46]\);
    
    \loop_all_sample.7.loop_all_chanel.1.sample_in_buf[118]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_693[118]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[118]\);
    
    \chanel_more.all_chanel.5.all_bit.3.sample_out_s2[68]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[50]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[68]\);
    
    \loop_all_sample.11.loop_all_chanel.5.sample_in_buf_RNO[42]\ : 
        MX2
      port map(A => \sample_in_buf[24]\, B => sample_5(11), S => 
        sample_val_delay, Y => \sample_in_buf_405[42]\);
    
    \chanel_more.all_chanel.3.all_bit.12.sample_out_s2[95]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[77]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[95]\);
    
    \loop_all_sample.1.loop_all_chanel.0.sample_in_buf_RNO[142]\ : 
        MX2
      port map(A => \sample_in_buf[124]\, B => sample_0(1), S => 
        sample_val_delay, Y => \sample_in_buf_1085[142]\);
    
    \loop_all_sample.12.loop_all_chanel.6.sample_in_buf[23]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_333[23]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[23]\);
    
    \chanel_more.all_chanel.5.all_bit.15.sample_out_s2[56]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[38]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[56]\);
    
    \loop_all_sample.4.loop_all_chanel.0.sample_in_buf[139]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_893[139]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[139]\);
    
    \chanel_more.all_chanel.6.all_bit.5.sample_out_s2[48]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[30]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[48]\);
    
    \loop_all_sample.4.loop_all_chanel.4.sample_in_buf[67]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_861[67]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[67]\);
    
    \loop_all_sample.12.loop_all_chanel.0.sample_in_buf_RNO[131]\ : 
        MX2
      port map(A => \sample_in_buf[113]\, B => sample_0(12), S
         => sample_val_delay, Y => \sample_in_buf_381[131]\);
    
    \chanel_more.all_chanel.4.all_bit.2.sample_out_s2[87]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[69]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[87]\);
    
    \loop_all_sample.5.loop_all_chanel.0.sample_in_buf_RNO[138]\ : 
        MX2
      port map(A => \sample_in_buf[120]\, B => sample_0(5), S => 
        sample_val_delay, Y => \sample_in_buf_829[138]\);
    
    \chanel_more.all_chanel.7.all_bit.5.sample_out_s2[30]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[12]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[30]\);
    
    \chanel_more.all_chanel.5.all_bit.14.sample_out_s2[57]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[39]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[57]\);
    
    \loop_all_sample.9.loop_all_chanel.5.sample_in_buf_RNO[44]\ : 
        MX2
      port map(A => \sample_in_buf[26]\, B => sample_5(9), S => 
        sample_val_delay, Y => \sample_in_buf_533[44]\);
    
    \chanel_more.all_chanel.3.all_bit.2.sample_out_s2[105]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[87]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[105]\);
    
    \loop_all_sample.5.loop_all_chanel.2.sample_in_buf[102]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_813[102]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[102]\);
    
    \chanel_HIGH.10.sample_out_s2[7]\ : DFN1E1C0
      port map(D => \sample_out_s[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[7]\);
    
    \chanel_more.all_chanel.6.all_bit.13.sample_out_s2[40]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[22]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[40]\);
    
    \chanel_more.all_chanel.5.all_bit.12.sample_out_s2[59]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[41]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[59]\);
    
    \loop_all_sample.14.loop_all_chanel.3.sample_in_buf[75]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_229[75]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[75]\);
    
    \loop_all_sample.14.loop_all_chanel.2.sample_in_buf_RNO[93]\ : 
        MX2
      port map(A => \sample_in_buf[75]\, B => sample_2(14), S => 
        sample_val_delay, Y => \sample_in_buf_237[93]\);
    
    \loop_all_sample.10.loop_all_chanel.5.sample_in_buf_RNO[43]\ : 
        MX2
      port map(A => \sample_in_buf[25]\, B => sample_5(10), S => 
        sample_val_delay, Y => \sample_in_buf_469[43]\);
    
    \loop_all_sample.0.loop_all_chanel.7.sample_in_buf[17]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1093[17]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[17]\);
    
    \loop_all_sample.6.loop_all_chanel.3.sample_in_buf_RNO[83]\ : 
        MX2
      port map(A => \sample_in_buf[65]\, B => sample_3(6), S => 
        sample_val_delay, Y => \sample_in_buf_741[83]\);
    
    \loop_all_sample.5.loop_all_chanel.6.sample_in_buf[30]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_781[30]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[30]\);
    
    \loop_all_sample.13.loop_all_chanel.0.sample_in_buf[130]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_317[130]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[130]\);
    
    \loop_all_sample.10.loop_all_chanel.7.sample_in_buf[7]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_453[7]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[7]\);
    
    \loop_all_sample.0.loop_all_chanel.0.sample_in_buf_RNO[143]\ : 
        MX2
      port map(A => \sample_in_buf[125]\, B => sample_0(0), S => 
        sample_val_delay, Y => \sample_in_buf_1149[143]\);
    
    \chanel_more.all_chanel.4.all_bit.12.sample_out_s2[77]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[59]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[77]\);
    
    \loop_all_sample.2.loop_all_chanel.6.sample_in_buf_RNO[33]\ : 
        MX2
      port map(A => \sample_in_buf[15]\, B => sample_6(2), S => 
        sample_val_delay, Y => \sample_in_buf_973[33]\);
    
    \chanel_more.all_chanel.5.all_bit.5.sample_out_s2[66]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[48]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[66]\);
    
    \loop_all_sample.6.loop_all_chanel.1.sample_in_buf[119]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_757[119]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[119]\);
    
    \loop_all_sample.0.loop_all_chanel.5.sample_in_buf[53]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1109[53]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[53]\);
    
    \loop_all_sample.17.loop_all_chanel.6.sample_in_buf_RNO[18]\ : 
        MX2
      port map(A => \sample_in_buf[0]\, B => sample_6(15), S => 
        sample_val_delay, Y => \sample_in_buf_13[18]\);
    
    \chanel_more.all_chanel.6.all_bit.4.sample_out_s2[49]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[31]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[49]\);
    
    \chanel_more.all_chanel.5.all_bit.1.sample_out_s2[70]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[52]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[70]\);
    
    \loop_all_sample.17.loop_all_chanel.7.sample_in_buf[0]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[0]\);
    
    \chanel_more.all_chanel.1.all_bit.14.sample_out_s2[129]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[111]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_127);
    
    \loop_all_sample.5.loop_all_chanel.1.sample_in_buf_RNO[120]\ : 
        MX2
      port map(A => \sample_in_buf[102]\, B => sample_1(5), S => 
        sample_val_delay, Y => \sample_in_buf_821[120]\);
    
    \loop_all_sample.0.loop_all_chanel.7.sample_in_buf_RNO[17]\ : 
        MX2
      port map(A => \sample_in_buf[143]\, B => sample_7(0), S => 
        sample_val_delay, Y => \sample_in_buf_1093[17]\);
    
    \loop_all_sample.12.loop_all_chanel.7.sample_in_buf[5]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_325[5]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[5]\);
    
    \chanel_more.all_chanel.3.all_bit.8.sample_out_s2[99]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[81]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[99]\);
    
    \chanel_more.all_chanel.4.all_bit.7.sample_out_s2[82]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[64]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[82]\);
    
    \loop_all_sample.10.loop_all_chanel.0.sample_in_buf[133]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_509[133]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[133]\);
    
    \loop_all_sample.3.loop_all_chanel.7.sample_in_buf[14]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_901[14]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[14]\);
    
    \chanel_HIGH.8.sample_out_s2[9]\ : DFN1E1C0
      port map(D => \sample_out_s[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[9]\);
    
    \chanel_more.all_chanel.5.all_bit.2.sample_out_s2[69]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[51]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[69]\);
    
    \chanel_more.all_chanel.1.all_bit.0.sample_out_s2[143]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[125]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_141);
    
    \chanel_more.all_chanel.1.all_bit.12.sample_out_s2[131]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[113]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_129);
    
    \chanel_HIGH.3.sample_out_s2[14]\ : DFN1E1C0
      port map(D => \sample_out_s[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[14]\);
    
    \chanel_more.all_chanel.7.all_bit.12.sample_out_s2[23]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[5]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[23]\);
    
    \loop_all_sample.8.loop_all_chanel.1.sample_in_buf_RNO[117]\ : 
        MX2
      port map(A => \sample_in_buf[99]\, B => sample_1(8), S => 
        sample_val_delay, Y => \sample_in_buf_629[117]\);
    
    \loop_all_sample.10.loop_all_chanel.0.sample_in_buf_RNO[133]\ : 
        MX2
      port map(A => \sample_in_buf[115]\, B => sample_0(10), S
         => sample_val_delay, Y => \sample_in_buf_509[133]\);
    
    \loop_all_sample.11.loop_all_chanel.3.sample_in_buf[78]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_421[78]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[78]\);
    
    \chanel_HIGH.11.sample_out_s2[6]\ : DFN1E1C0
      port map(D => \sample_out_s[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_out_rot_s_0, Q => 
        \sample_filter_v2_out[6]\);
    
    \loop_all_sample.10.loop_all_chanel.3.sample_in_buf_RNO[79]\ : 
        MX2
      port map(A => \sample_in_buf[61]\, B => sample_3(10), S => 
        sample_val_delay, Y => \sample_in_buf_485[79]\);
    
    \chanel_more.all_chanel.1.all_bit.11.sample_out_s2[132]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[114]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_130);
    
    \chanel_more.all_chanel.1.all_bit.10.sample_out_s2[133]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[115]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_0, Q => 
        sample_filter_v2_out_131);
    
    \loop_all_sample.13.loop_all_chanel.1.sample_in_buf_RNO[112]\ : 
        MX2
      port map(A => \sample_in_buf[94]\, B => sample_1(13), S => 
        sample_val_delay, Y => \sample_in_buf_309[112]\);
    
    \loop_all_sample.6.loop_all_chanel.3.sample_in_buf[83]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_741[83]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[83]\);
    
    \loop_all_sample.2.loop_all_chanel.3.sample_in_buf_RNO[87]\ : 
        MX2
      port map(A => \sample_in_buf[69]\, B => sample_3(2), S => 
        sample_val_delay, Y => \sample_in_buf_997[87]\);
    
    \loop_all_sample.1.loop_all_chanel.5.sample_in_buf[52]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_1045[52]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[52]\);
    
    \chanel_more.all_chanel.7.all_bit.0.sample_out_s2[35]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[17]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[35]\);
    
    \chanel_more.all_chanel.4.all_bit.14.sample_out_s2[75]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[57]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[75]\);
    
    \chanel_more.all_chanel.2.all_bit.4.sample_out_s2[121]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[103]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[121]\);
    
    \chanel_more.all_chanel.2.all_bit.12.sample_out_s2[113]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[95]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        \sample_filter_v2_out[113]\);
    
    \chanel_more.all_chanel.1.all_bit.7.sample_out_s2[136]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[118]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_134);
    
    \chanel_more.all_chanel.1.all_bit.2.sample_out_s2[141]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[123]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_1, Q => 
        sample_filter_v2_out_139);
    
    \loop_all_sample.6.loop_all_chanel.2.sample_in_buf_RNO[101]\ : 
        MX2
      port map(A => \sample_in_buf[83]\, B => sample_2(6), S => 
        sample_val_delay, Y => \sample_in_buf_749[101]\);
    
    \chanel_more.all_chanel.5.all_bit.11.sample_out_s2[60]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[42]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_3, Q => 
        \sample_filter_v2_out[60]\);
    
    \loop_all_sample.1.loop_all_chanel.1.sample_in_buf_RNO[124]\ : 
        MX2
      port map(A => \sample_in_buf[106]\, B => sample_1(1), S => 
        sample_val_delay, Y => \sample_in_buf_1077[124]\);
    
    IIR_CEL_CTRLR_v2_CONTROL_1 : IIR_CEL_CTRLR_v2_CONTROL
      port map(alu_ctrl(2) => \alu_ctrl[2]\, alu_ctrl(1) => 
        \alu_ctrl[1]\, alu_ctrl(0) => \alu_ctrl[0]\, 
        ram_sel_Wdata(1) => \ram_sel_Wdata[1]\, ram_sel_Wdata(0)
         => \ram_sel_Wdata[0]\, waddr_previous(1) => 
        \waddr_previous[1]\, waddr_previous(0) => 
        \waddr_previous[0]\, in_sel_src(1) => \in_sel_src[1]\, 
        in_sel_src(0) => \in_sel_src[0]\, S_i_0(33) => 
        \S_i_0[33]\, S(8) => \S[8]\, alu_sel_coeff(4) => 
        \alu_sel_coeff[4]\, alu_sel_coeff(3) => 
        \alu_sel_coeff[3]\, alu_sel_coeff(2) => 
        \alu_sel_coeff[2]\, alu_sel_coeff(1) => 
        \alu_sel_coeff[1]\, alu_sel_coeff(0) => 
        \alu_sel_coeff[0]\, alu_sel_coeff_0_2 => 
        \alu_sel_coeff_0[2]\, alu_sel_coeff_0_0 => 
        \alu_sel_coeff_0[0]\, sample_out_rot_s => 
        sample_out_rot_s, sample_out_val_s => sample_out_val_s, 
        raddr_rst => raddr_rst, alu_sel_input => alu_sel_input, 
        raddr_add1 => raddr_add1, sample_val_delay => 
        sample_val_delay, ram_write => ram_write, ram_write_i => 
        ram_write_i, un1_sample_in_rotate => un1_sample_in_rotate, 
        sample_out_rot_s_0 => sample_out_rot_s_0, 
        sample_out_rot_s_1 => sample_out_rot_s_1, 
        sample_out_rot_s_2 => sample_out_rot_s_2, 
        sample_out_rot_s_3 => sample_out_rot_s_3, 
        sample_out_rot_s_4 => sample_out_rot_s_4, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    \loop_all_sample.7.loop_all_chanel.3.sample_in_buf_RNO[82]\ : 
        MX2
      port map(A => \sample_in_buf[64]\, B => sample_3(7), S => 
        sample_val_delay, Y => \sample_in_buf_677[82]\);
    
    \chanel_more.all_chanel.7.all_bit.8.sample_out_s2[27]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[9]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[27]\);
    
    \chanel_more.all_chanel.6.all_bit.7.sample_out_s2[46]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[28]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_4, Q => 
        \sample_filter_v2_out[46]\);
    
    \loop_all_sample.7.loop_all_chanel.3.sample_in_buf[82]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_677[82]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[82]\);
    
    \loop_all_sample.17.loop_all_chanel.0.sample_in_buf[126]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_61[126]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[128]\);
    
    \loop_all_sample.11.loop_all_chanel.4.sample_in_buf[60]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_413[60]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[60]\);
    
    \loop_all_sample.3.loop_all_chanel.6.sample_in_buf_RNO[32]\ : 
        MX2
      port map(A => \sample_in_buf[14]\, B => sample_6(3), S => 
        sample_val_delay, Y => \sample_in_buf_909[32]\);
    
    \loop_all_sample.17.loop_all_chanel.1.sample_in_buf_RNO[108]\ : 
        MX2
      port map(A => \sample_in_buf[90]\, B => sample_1(15), S => 
        sample_val_delay, Y => \sample_in_buf_53[108]\);
    
    \loop_all_sample.8.loop_all_chanel.6.sample_in_buf_RNO[27]\ : 
        MX2
      port map(A => \sample_in_buf[9]\, B => sample_6(8), S => 
        sample_val_delay, Y => \sample_in_buf_589[27]\);
    
    \loop_all_sample.5.loop_all_chanel.4.sample_in_buf[66]\ : 
        DFN1E1C0
      port map(D => \sample_in_buf_797[66]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => un1_sample_in_rotate, Q => 
        \sample_in_buf[66]\);
    
    \loop_all_sample.14.loop_all_chanel.1.sample_in_buf_RNO[111]\ : 
        MX2
      port map(A => \sample_in_buf[93]\, B => sample_1(14), S => 
        sample_val_delay, Y => \sample_in_buf_245[111]\);
    
    \chanel_more.all_chanel.2.all_bit.8.sample_out_s2[117]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[99]\, CLK => HCLK_c, 
        CLR => HRESETn_c, E => sample_out_rot_s_2, Q => 
        \sample_filter_v2_out[117]\);
    
    \chanel_more.all_chanel.7.all_bit.11.sample_out_s2[24]\ : 
        DFN1E1C0
      port map(D => \sample_filter_v2_out[6]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sample_out_rot_s, Q => 
        \sample_filter_v2_out[24]\);
    
    \loop_all_sample.8.loop_all_chanel.2.sample_in_buf_RNO[99]\ : 
        MX2
      port map(A => \sample_in_buf[81]\, B => sample_2(8), S => 
        sample_val_delay, Y => \sample_in_buf_621[99]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Downsampling_6_16_256 is

    port( sample_f1          : in    std_logic_vector(111 downto 80);
          sample_f1_wdata_95 : in    std_logic;
          sample_f1_wdata_94 : in    std_logic;
          sample_f1_wdata_93 : in    std_logic;
          sample_f1_wdata_92 : in    std_logic;
          sample_f1_wdata_91 : in    std_logic;
          sample_f1_wdata_90 : in    std_logic;
          sample_f1_wdata_89 : in    std_logic;
          sample_f1_wdata_88 : in    std_logic;
          sample_f1_wdata_87 : in    std_logic;
          sample_f1_wdata_86 : in    std_logic;
          sample_f1_wdata_85 : in    std_logic;
          sample_f1_wdata_84 : in    std_logic;
          sample_f1_wdata_83 : in    std_logic;
          sample_f1_wdata_82 : in    std_logic;
          sample_f1_wdata_81 : in    std_logic;
          sample_f1_wdata_80 : in    std_logic;
          sample_f1_wdata_79 : in    std_logic;
          sample_f1_wdata_78 : in    std_logic;
          sample_f1_wdata_77 : in    std_logic;
          sample_f1_wdata_76 : in    std_logic;
          sample_f1_wdata_75 : in    std_logic;
          sample_f1_wdata_74 : in    std_logic;
          sample_f1_wdata_73 : in    std_logic;
          sample_f1_wdata_72 : in    std_logic;
          sample_f1_wdata_71 : in    std_logic;
          sample_f1_wdata_70 : in    std_logic;
          sample_f1_wdata_69 : in    std_logic;
          sample_f1_wdata_68 : in    std_logic;
          sample_f1_wdata_67 : in    std_logic;
          sample_f1_wdata_66 : in    std_logic;
          sample_f1_wdata_65 : in    std_logic;
          sample_f1_wdata_64 : in    std_logic;
          sample_f1_wdata_63 : in    std_logic;
          sample_f1_wdata_62 : in    std_logic;
          sample_f1_wdata_61 : in    std_logic;
          sample_f1_wdata_60 : in    std_logic;
          sample_f1_wdata_59 : in    std_logic;
          sample_f1_wdata_58 : in    std_logic;
          sample_f1_wdata_57 : in    std_logic;
          sample_f1_wdata_56 : in    std_logic;
          sample_f1_wdata_55 : in    std_logic;
          sample_f1_wdata_54 : in    std_logic;
          sample_f1_wdata_53 : in    std_logic;
          sample_f1_wdata_52 : in    std_logic;
          sample_f1_wdata_51 : in    std_logic;
          sample_f1_wdata_50 : in    std_logic;
          sample_f1_wdata_49 : in    std_logic;
          sample_f1_wdata_48 : in    std_logic;
          sample_f1_wdata_15 : in    std_logic;
          sample_f1_wdata_14 : in    std_logic;
          sample_f1_wdata_13 : in    std_logic;
          sample_f1_wdata_12 : in    std_logic;
          sample_f1_wdata_11 : in    std_logic;
          sample_f1_wdata_10 : in    std_logic;
          sample_f1_wdata_9  : in    std_logic;
          sample_f1_wdata_8  : in    std_logic;
          sample_f1_wdata_7  : in    std_logic;
          sample_f1_wdata_6  : in    std_logic;
          sample_f1_wdata_5  : in    std_logic;
          sample_f1_wdata_4  : in    std_logic;
          sample_f1_wdata_3  : in    std_logic;
          sample_f1_wdata_2  : in    std_logic;
          sample_f1_wdata_1  : in    std_logic;
          sample_f1_wdata_0  : in    std_logic;
          sample_f3_wdata    : out   std_logic_vector(95 downto 0);
          sample_f1_val      : in    std_logic;
          HCLK_c             : in    std_logic;
          sample_f3_val      : out   std_logic;
          HRESETn_c          : in    std_logic;
          sample_f1_val_0    : in    std_logic
        );

end Downsampling_6_16_256;

architecture DEF_ARCH of Downsampling_6_16_256 is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un2_sample_in_val_0, un2_sample_in_val_23, 
        un2_sample_in_val_22, un2_sample_in_val_24, 
        sample_out_0_sqmuxa_2, sample_out_0_sqmuxa_1, 
        sample_out_0_sqmuxa_0, N_137, \counter[1]_net_1\, 
        \counter[0]_net_1\, N_129, \counter[3]_net_1\, 
        \DWACT_FDEC_E[0]\, N_106, \counter[8]_net_1\, 
        \DWACT_FDEC_E[4]\, N_91, \DWACT_FDEC_E[7]\, 
        \DWACT_FDEC_E[6]\, un2_sample_in_val_15, 
        un2_sample_in_val_14, un2_sample_in_val_20, 
        un2_sample_in_val_9, un2_sample_in_val_8, 
        un2_sample_in_val_19, un2_sample_in_val_5, 
        un2_sample_in_val_4, un2_sample_in_val_17, 
        un2_sample_in_val_13, \counter[24]_net_1\, 
        un2_sample_in_val_11, \counter[15]_net_1\, 
        \counter[12]_net_1\, un2_sample_in_val_7, 
        \counter[22]_net_1\, \counter[19]_net_1\, 
        un2_sample_in_val_3, \counter[23]_net_1\, 
        \counter[20]_net_1\, un2_sample_in_val_1, 
        \counter[11]_net_1\, \counter[27]_net_1\, 
        \counter[18]_net_1\, \counter[21]_net_1\, 
        \counter[9]_net_1\, \counter[4]_net_1\, 
        \counter[6]_net_1\, \counter[25]_net_1\, 
        \counter[2]_net_1\, \counter[13]_net_1\, 
        \counter[16]_net_1\, \counter[7]_net_1\, 
        \counter[10]_net_1\, \counter[26]_net_1\, 
        \counter[5]_net_1\, \counter[14]_net_1\, 
        \counter[17]_net_1\, un2_sample_in_val, 
        sample_out_0_sqmuxa, \counter_4[8]\, I_45_2, 
        \counter_4[9]\, I_52_2, \counter_4[10]\, I_56_2, 
        \counter_4[11]\, I_66_2, \counter_4[12]\, I_73_2, 
        \counter_4[13]\, I_77_2, \counter_4[14]\, I_84_2, 
        \counter_4[15]\, I_91_2, \counter_4[16]\, I_98_2, 
        \counter_4[17]\, I_105_2, \counter_4[18]\, I_115_2, 
        \counter_4[19]\, I_122_2, \counter_4[20]\, I_129_2, 
        \counter_4[21]\, I_136_2, \counter_4[22]\, I_143_2, 
        \counter_4[23]\, I_156_2, \counter_4[24]\, I_166_2, 
        \counter_4[25]\, I_173_2, \counter_4[26]\, I_186_2, 
        \counter_4[27]\, I_196_2, sample_out_val_4, I_4_2, I_5_2, 
        I_9_2, I_13_2, I_20_2, I_24_2, I_31_3, I_38_2, N_4, 
        \DWACT_FDEC_E[29]\, \DWACT_FDEC_E[30]\, 
        \DWACT_FDEC_E[23]\, \DWACT_FDEC_E[15]\, 
        \DWACT_FDEC_E[17]\, \DWACT_FDEC_E[22]\, N_11, 
        \DWACT_FDEC_E[21]\, \DWACT_FDEC_E[9]\, \DWACT_FDEC_E[12]\, 
        \DWACT_FDEC_E[20]\, N_20, \DWACT_FDEC_E[13]\, 
        \DWACT_FDEC_E[19]\, N_25, \DWACT_FDEC_E[18]\, N_32, 
        \DWACT_FDEC_E[33]\, \DWACT_FDEC_E[34]\, \DWACT_FDEC_E[2]\, 
        \DWACT_FDEC_E[5]\, N_41, \DWACT_FDEC_E[28]\, 
        \DWACT_FDEC_E[16]\, N_46, N_51, \DWACT_FDEC_E[14]\, N_56, 
        N_61, \DWACT_FDEC_E[10]\, N_68, \DWACT_FDEC_E[11]\, N_73, 
        N_78, N_83, \DWACT_FDEC_E[8]\, N_88, N_96, N_103, 
        \DWACT_FDEC_E[3]\, N_111, N_116, N_121, \DWACT_FDEC_E[1]\, 
        N_126, N_134, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \counter[19]\ : DFN1E1C0
      port map(D => \counter_4[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[19]_net_1\);
    
    \counter_RNI8DTE[12]\ : NOR3C
      port map(A => un2_sample_in_val_9, B => un2_sample_in_val_8, 
        C => un2_sample_in_val_19, Y => un2_sample_in_val_23);
    
    \sample_out[22]\ : DFN1E1
      port map(D => sample_f1_wdata_73, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(73));
    
    \sample_out[20]\ : DFN1E1
      port map(D => sample_f1_wdata_75, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(75));
    
    \sample_out[13]\ : DFN1E1
      port map(D => sample_f1_wdata_82, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(82));
    
    \sample_out[1]\ : DFN1E1
      port map(D => sample_f1_wdata_94, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(94));
    
    \sample_out[19]\ : DFN1E1
      port map(D => sample_f1_wdata_76, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(76));
    
    un3_counter_I_142 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[16]\, Y => N_41);
    
    \sample_out[61]\ : DFN1E1
      port map(D => sample_f1(93), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(34));
    
    \sample_out[66]\ : DFN1E1
      port map(D => sample_f1(98), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(29));
    
    \sample_out[73]\ : DFN1E1
      port map(D => sample_f1(105), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(22));
    
    \sample_out[79]\ : DFN1E1
      port map(D => sample_f1(111), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(16));
    
    \sample_out[38]\ : DFN1E1
      port map(D => sample_f1_wdata_57, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(57));
    
    un3_counter_I_27 : OR2
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        Y => \DWACT_FDEC_E[1]\);
    
    \sample_out[95]\ : DFN1E1
      port map(D => sample_f1_wdata_0, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(0));
    
    \counter_RNO[11]\ : NOR2B
      port map(A => I_66_2, B => un2_sample_in_val_0, Y => 
        \counter_4[11]\);
    
    \sample_out[34]\ : DFN1E1
      port map(D => sample_f1_wdata_61, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(61));
    
    un3_counter_I_4 : INV
      port map(A => \counter[0]_net_1\, Y => I_4_2);
    
    \counter[11]\ : DFN1E1C0
      port map(D => \counter_4[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[11]_net_1\);
    
    un3_counter_I_94 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, Y
         => \DWACT_FDEC_E[10]\);
    
    un3_counter_I_186 : XNOR2
      port map(A => N_11, B => \counter[26]_net_1\, Y => I_186_2);
    
    \counter_RNO[15]\ : NOR2B
      port map(A => I_91_2, B => un2_sample_in_val_0, Y => 
        \counter_4[15]\);
    
    un3_counter_I_108 : OR3
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        C => \counter[17]_net_1\, Y => \DWACT_FDEC_E[12]\);
    
    un3_counter_I_121 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \counter[18]_net_1\, Y => N_56);
    
    \sample_out[51]\ : DFN1E1
      port map(D => sample_f1(83), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(44));
    
    \sample_out[56]\ : DFN1E1
      port map(D => sample_f1(88), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(39));
    
    un3_counter_I_176 : OR2
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        Y => \DWACT_FDEC_E[20]\);
    
    \sample_out[0]\ : DFN1E1
      port map(D => sample_f1_wdata_95, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(95));
    
    \counter[6]\ : DFN1E1C0
      port map(D => I_31_3, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f1_val, Q => \counter[6]_net_1\);
    
    un3_counter_I_48 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => \DWACT_FDEC_E[4]\);
    
    un3_counter_I_114 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[10]\, 
        C => \DWACT_FDEC_E[12]\, Y => N_61);
    
    \counter[21]\ : DFN1E1C0
      port map(D => \counter_4[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[21]_net_1\);
    
    un3_counter_I_13 : XNOR2
      port map(A => N_134, B => \counter[3]_net_1\, Y => I_13_2);
    
    \sample_out[81]\ : DFN1E1
      port map(D => sample_f1_wdata_14, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(14));
    
    \sample_out[86]\ : DFN1E1
      port map(D => sample_f1_wdata_9, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(9));
    
    \counter[3]\ : DFN1E1C0
      port map(D => I_13_2, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f1_val, Q => \counter[3]_net_1\);
    
    \counter[2]\ : DFN1E1C0
      port map(D => I_9_2, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f1_val, Q => \counter[2]_net_1\);
    
    un3_counter_I_73 : XNOR2
      port map(A => N_91, B => \counter[12]_net_1\, Y => I_73_2);
    
    \counter_RNO[8]\ : NOR2B
      port map(A => I_45_2, B => un2_sample_in_val_0, Y => 
        \counter_4[8]\);
    
    \counter_RNO[13]\ : NOR2B
      port map(A => I_77_2, B => un2_sample_in_val_0, Y => 
        \counter_4[13]\);
    
    un3_counter_I_52 : XNOR2
      port map(A => N_106, B => \counter[9]_net_1\, Y => I_52_2);
    
    \sample_out[12]\ : DFN1E1
      port map(D => sample_f1_wdata_83, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(83));
    
    \sample_out[10]\ : DFN1E1
      port map(D => sample_f1_wdata_85, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(85));
    
    \sample_out[45]\ : DFN1E1
      port map(D => sample_f1_wdata_50, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(50));
    
    \counter_RNO[12]\ : NOR2B
      port map(A => I_73_2, B => un2_sample_in_val_0, Y => 
        \counter_4[12]\);
    
    \sample_out[72]\ : DFN1E1
      port map(D => sample_f1(104), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(23));
    
    \sample_out[33]\ : DFN1E1
      port map(D => sample_f1_wdata_62, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(62));
    
    \sample_out[39]\ : DFN1E1
      port map(D => sample_f1_wdata_56, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(56));
    
    \counter[17]\ : DFN1E1C0
      port map(D => \counter_4[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[17]_net_1\);
    
    \sample_out[70]\ : DFN1E1
      port map(D => sample_f1(102), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(25));
    
    un3_counter_I_41 : OR2
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        Y => \DWACT_FDEC_E[3]\);
    
    un3_counter_I_159 : OR3
      port map(A => \counter[21]_net_1\, B => \counter[22]_net_1\, 
        C => \counter[23]_net_1\, Y => \DWACT_FDEC_E[17]\);
    
    \counter[4]\ : DFN1E1C0
      port map(D => I_20_2, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f1_val, Q => \counter[4]_net_1\);
    
    un3_counter_I_5 : XNOR2
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        Y => I_5_2);
    
    un3_counter_I_125 : OR2
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        Y => \DWACT_FDEC_E[14]\);
    
    \counter[10]\ : DFN1E1C0
      port map(D => \counter_4[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[10]_net_1\);
    
    \sample_out[5]\ : DFN1E1
      port map(D => sample_f1_wdata_90, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(90));
    
    \sample_out[47]\ : DFN1E1
      port map(D => sample_f1_wdata_48, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(48));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter[13]\ : DFN1E1C0
      port map(D => \counter_4[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[13]_net_1\);
    
    un3_counter_I_62 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[6]\);
    
    \counter_RNIPKE[13]\ : NOR2
      port map(A => \counter[13]_net_1\, B => \counter[16]_net_1\, 
        Y => un2_sample_in_val_5);
    
    \sample_out[65]\ : DFN1E1
      port map(D => sample_f1(97), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(30));
    
    \counter_RNIBJN3[26]\ : NOR2
      port map(A => \counter[26]_net_1\, B => \counter[5]_net_1\, 
        Y => un2_sample_in_val_3);
    
    un3_counter_I_139 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        Y => \DWACT_FDEC_E[16]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sample_out[21]\ : DFN1E1
      port map(D => sample_f1_wdata_74, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(74));
    
    \counter[12]\ : DFN1E1C0
      port map(D => \counter_4[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[12]_net_1\);
    
    \sample_out[26]\ : DFN1E1
      port map(D => sample_f1_wdata_69, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(69));
    
    \sample_out[2]\ : DFN1E1
      port map(D => sample_f1_wdata_93, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(93));
    
    \counter[27]\ : DFN1E1C0
      port map(D => \counter_4[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[27]_net_1\);
    
    \counter_RNI2SB8[10]\ : NOR3C
      port map(A => un2_sample_in_val_5, B => un2_sample_in_val_4, 
        C => un2_sample_in_val_17, Y => un2_sample_in_val_22);
    
    un3_counter_I_111 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[28]\);
    
    \sample_out[67]\ : DFN1E1
      port map(D => sample_f1(99), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(28));
    
    \counter[20]\ : DFN1E1C0
      port map(D => \counter_4[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[20]_net_1\);
    
    \sample_out[94]\ : DFN1E1
      port map(D => sample_f1_wdata_1, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(1));
    
    un3_counter_I_166 : XNOR2
      port map(A => N_25, B => \counter[24]_net_1\, Y => I_166_2);
    
    \counter_RNO[17]\ : NOR2B
      port map(A => I_105_2, B => un2_sample_in_val, Y => 
        \counter_4[17]\);
    
    \counter[23]\ : DFN1E1C0
      port map(D => \counter_4[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[23]_net_1\);
    
    un3_counter_I_149 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[34]\);
    
    \sample_out[55]\ : DFN1E1
      port map(D => sample_f1(87), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(40));
    
    \counter[22]\ : DFN1E1C0
      port map(D => \counter_4[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[22]_net_1\);
    
    \counter[15]\ : DFN1E1C0
      port map(D => \counter_4[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[15]_net_1\);
    
    un3_counter_I_8 : OR2
      port map(A => \counter[1]_net_1\, B => \counter[0]_net_1\, 
        Y => N_137);
    
    un3_counter_I_185 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[21]\, Y => N_11);
    
    \counter_RNIH507[3]\ : NOR2
      port map(A => \counter[3]_net_1\, B => \counter[0]_net_1\, 
        Y => un2_sample_in_val_13);
    
    un3_counter_I_196 : XNOR2
      port map(A => N_4, B => \counter[27]_net_1\, Y => I_196_2);
    
    \sample_out[32]\ : DFN1E1
      port map(D => sample_f1_wdata_63, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(63));
    
    un3_counter_I_51 : OR2
      port map(A => \counter[8]_net_1\, B => \DWACT_FDEC_E[4]\, Y
         => N_106);
    
    un3_counter_I_122 : XNOR2
      port map(A => N_56, B => \counter[19]_net_1\, Y => I_122_2);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sample_out[57]\ : DFN1E1
      port map(D => sample_f1(89), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(38));
    
    \sample_out[30]\ : DFN1E1
      port map(D => sample_f1_wdata_65, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(65));
    
    \counter_RNO[14]\ : NOR2B
      port map(A => I_84_2, B => un2_sample_in_val_0, Y => 
        \counter_4[14]\);
    
    \sample_out[85]\ : DFN1E1
      port map(D => sample_f1_wdata_10, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(10));
    
    \counter_RNIO507[4]\ : NOR2
      port map(A => \counter[4]_net_1\, B => \counter[6]_net_1\, 
        Y => un2_sample_in_val_8);
    
    \counter[1]\ : DFN1E1C0
      port map(D => I_5_2, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f1_val, Q => \counter[1]_net_1\);
    
    \counter_RNO[26]\ : NOR2B
      port map(A => I_186_2, B => un2_sample_in_val, Y => 
        \counter_4[26]\);
    
    \sample_out[4]\ : DFN1E1
      port map(D => sample_f1_wdata_91, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(91));
    
    \counter_RNI0MBF1_2[10]\ : NOR3B
      port map(A => sample_f1_val_0, B => HRESETn_c, C => 
        un2_sample_in_val_0, Y => sample_out_0_sqmuxa_1);
    
    \counter[25]\ : DFN1E1C0
      port map(D => \counter_4[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[25]_net_1\);
    
    sample_out_val : DFN1C0
      port map(D => sample_out_val_4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f3_val);
    
    \sample_out[87]\ : DFN1E1
      port map(D => sample_f1_wdata_8, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(8));
    
    un3_counter_I_115 : XNOR2
      port map(A => N_61, B => \counter[18]_net_1\, Y => I_115_2);
    
    un3_counter_I_87 : OR3
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        C => \counter[14]_net_1\, Y => \DWACT_FDEC_E[9]\);
    
    un3_counter_I_173 : XNOR2
      port map(A => N_20, B => \counter[25]_net_1\, Y => I_173_2);
    
    \sample_out[48]\ : DFN1E1
      port map(D => sample_f1(80), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(47));
    
    un3_counter_I_38 : XNOR2
      port map(A => N_116, B => \counter[7]_net_1\, Y => I_38_2);
    
    \sample_out[93]\ : DFN1E1
      port map(D => sample_f1_wdata_2, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(2));
    
    \sample_out[11]\ : DFN1E1
      port map(D => sample_f1_wdata_84, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(84));
    
    \sample_out[16]\ : DFN1E1
      port map(D => sample_f1_wdata_79, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(79));
    
    \counter[5]\ : DFN1E1C0
      port map(D => I_24_2, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f1_val, Q => \counter[5]_net_1\);
    
    \sample_out[44]\ : DFN1E1
      port map(D => sample_f1_wdata_51, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(51));
    
    \sample_out[71]\ : DFN1E1
      port map(D => sample_f1(103), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(24));
    
    \sample_out[76]\ : DFN1E1
      port map(D => sample_f1(108), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(19));
    
    un3_counter_I_37 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \counter[6]_net_1\, Y => N_116);
    
    \counter_RNO[10]\ : NOR2B
      port map(A => I_56_2, B => un2_sample_in_val_0, Y => 
        \counter_4[10]\);
    
    \counter_RNIRSE[14]\ : NOR2
      port map(A => \counter[14]_net_1\, B => \counter[17]_net_1\, 
        Y => un2_sample_in_val_1);
    
    un3_counter_I_9 : XNOR2
      port map(A => N_137, B => \counter[2]_net_1\, Y => I_9_2);
    
    \counter_RNO[21]\ : NOR2B
      port map(A => I_136_2, B => un2_sample_in_val, Y => 
        \counter_4[21]\);
    
    un3_counter_I_20 : XNOR2
      port map(A => N_129, B => \counter[4]_net_1\, Y => I_20_2);
    
    un3_counter_I_182 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[30]\);
    
    \sample_out[68]\ : DFN1E1
      port map(D => sample_f1(100), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(27));
    
    \sample_out[25]\ : DFN1E1
      port map(D => sample_f1_wdata_70, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(70));
    
    un3_counter_I_56 : XNOR2
      port map(A => N_103, B => \counter[10]_net_1\, Y => I_56_2);
    
    \counter[16]\ : DFN1E1C0
      port map(D => \counter_4[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[16]_net_1\);
    
    \counter_RNO[25]\ : NOR2B
      port map(A => I_173_2, B => un2_sample_in_val, Y => 
        \counter_4[25]\);
    
    un3_counter_I_172 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[19]\, Y => N_20);
    
    un3_counter_I_104 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \DWACT_FDEC_E[11]\, Y => N_68);
    
    \sample_out[64]\ : DFN1E1
      port map(D => sample_f1(96), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(31));
    
    un3_counter_I_31 : XNOR2
      port map(A => N_121, B => \counter[6]_net_1\, Y => I_31_3);
    
    \counter_RNIH1T[12]\ : NOR3A
      port map(A => un2_sample_in_val_11, B => 
        \counter[15]_net_1\, C => \counter[12]_net_1\, Y => 
        un2_sample_in_val_19);
    
    \counter_RNI0G54[20]\ : NOR3A
      port map(A => un2_sample_in_val_3, B => \counter[23]_net_1\, 
        C => \counter[20]_net_1\, Y => un2_sample_in_val_15);
    
    un3_counter_I_98 : XNOR2
      port map(A => N_73, B => \counter[16]_net_1\, Y => I_98_2);
    
    un3_counter_I_23 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \counter[3]_net_1\, C
         => \counter[4]_net_1\, Y => N_126);
    
    \sample_out[27]\ : DFN1E1
      port map(D => sample_f1_wdata_68, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(68));
    
    un3_counter_I_59 : OR3
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        C => \counter[8]_net_1\, Y => \DWACT_FDEC_E[5]\);
    
    \counter_RNI6RM3[10]\ : NOR2
      port map(A => \counter[7]_net_1\, B => \counter[10]_net_1\, 
        Y => un2_sample_in_val_4);
    
    un3_counter_I_12 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => N_134);
    
    un3_counter_I_165 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[18]\, Y => N_25);
    
    un3_counter_I_156 : XNOR2
      port map(A => N_32, B => \counter[23]_net_1\, Y => I_156_2);
    
    un3_counter_I_97 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \counter[15]_net_1\, Y => N_73);
    
    un3_counter_I_128 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[14]\, Y => N_51);
    
    un3_counter_I_72 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[6]\, Y
         => N_91);
    
    \sample_out[58]\ : DFN1E1
      port map(D => sample_f1(90), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(37));
    
    \counter_RNI7FN3[25]\ : NOR2
      port map(A => \counter[25]_net_1\, B => \counter[2]_net_1\, 
        Y => un2_sample_in_val_7);
    
    \counter[26]\ : DFN1E1C0
      port map(D => \counter_4[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[26]_net_1\);
    
    un3_counter_I_66 : XNOR2
      port map(A => N_96, B => \counter[11]_net_1\, Y => I_66_2);
    
    \counter_RNO[23]\ : NOR2B
      port map(A => I_156_2, B => un2_sample_in_val, Y => 
        \counter_4[23]\);
    
    \sample_out[54]\ : DFN1E1
      port map(D => sample_f1(86), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(41));
    
    \sample_out[43]\ : DFN1E1
      port map(D => sample_f1_wdata_52, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(52));
    
    \sample_out[49]\ : DFN1E1
      port map(D => sample_f1(81), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(46));
    
    \counter_RNI0MBF1_0[10]\ : NOR3B
      port map(A => sample_f1_val_0, B => HRESETn_c, C => 
        un2_sample_in_val_0, Y => sample_out_0_sqmuxa_0);
    
    un3_counter_I_45 : XNOR2
      port map(A => N_111, B => \counter[8]_net_1\, Y => I_45_2);
    
    un3_counter_I_24 : XNOR2
      port map(A => N_126, B => \counter[5]_net_1\, Y => I_24_2);
    
    un3_counter_I_195 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[23]\, Y => N_4);
    
    \sample_out[92]\ : DFN1E1
      port map(D => sample_f1_wdata_3, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(3));
    
    \counter[14]\ : DFN1E1C0
      port map(D => \counter_4[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val_0, Q => \counter[14]_net_1\);
    
    un3_counter_I_136 : XNOR2
      port map(A => N_46, B => \counter[21]_net_1\, Y => I_136_2);
    
    \sample_out[88]\ : DFN1E1
      port map(D => sample_f1_wdata_7, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(7));
    
    \sample_out[90]\ : DFN1E1
      port map(D => sample_f1_wdata_5, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(5));
    
    un3_counter_I_91 : XNOR2
      port map(A => N_78, B => \counter[15]_net_1\, Y => I_91_2);
    
    \counter_RNO[22]\ : NOR2B
      port map(A => I_143_2, B => un2_sample_in_val, Y => 
        \counter_4[22]\);
    
    \sample_out[31]\ : DFN1E1
      port map(D => sample_f1_wdata_64, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(64));
    
    \sample_out[36]\ : DFN1E1
      port map(D => sample_f1_wdata_59, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(59));
    
    un3_counter_I_69 : OR3
      port map(A => \counter[9]_net_1\, B => \counter[10]_net_1\, 
        C => \counter[11]_net_1\, Y => \DWACT_FDEC_E[7]\);
    
    \sample_out[84]\ : DFN1E1
      port map(D => sample_f1_wdata_11, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(11));
    
    \sample_out[63]\ : DFN1E1
      port map(D => sample_f1(95), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(32));
    
    \sample_out[69]\ : DFN1E1
      port map(D => sample_f1(101), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(26));
    
    \sample_out[15]\ : DFN1E1
      port map(D => sample_f1_wdata_80, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(80));
    
    un3_counter_I_129 : XNOR2
      port map(A => N_51, B => \counter[20]_net_1\, Y => I_129_2);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un3_counter_I_146 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        C => \counter[22]_net_1\, Y => \DWACT_FDEC_E[33]\);
    
    \counter[24]\ : DFN1E1C0
      port map(D => \counter_4[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[24]_net_1\);
    
    un3_counter_I_101 : OR2
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        Y => \DWACT_FDEC_E[11]\);
    
    \sample_out[75]\ : DFN1E1
      port map(D => sample_f1(107), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(20));
    
    \counter_RNIMGNA[24]\ : NOR3A
      port map(A => un2_sample_in_val_13, B => \counter[1]_net_1\, 
        C => \counter[24]_net_1\, Y => un2_sample_in_val_20);
    
    un3_counter_I_162 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        Y => \DWACT_FDEC_E[18]\);
    
    \counter_RNIKN371[10]\ : OR3C
      port map(A => un2_sample_in_val_23, B => 
        un2_sample_in_val_22, C => un2_sample_in_val_24, Y => 
        un2_sample_in_val_0);
    
    un3_counter_I_77 : XNOR2
      port map(A => N_88, B => \counter[13]_net_1\, Y => I_77_2);
    
    \sample_out[17]\ : DFN1E1
      port map(D => sample_f1_wdata_78, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(78));
    
    \counter_RNO[18]\ : NOR2B
      port map(A => I_115_2, B => un2_sample_in_val, Y => 
        \counter_4[18]\);
    
    un3_counter_I_44 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => N_111);
    
    \sample_out[77]\ : DFN1E1
      port map(D => sample_f1(109), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(18));
    
    \counter_RNI0MBF1[10]\ : NOR3B
      port map(A => sample_f1_val_0, B => HRESETn_c, C => 
        un2_sample_in_val_0, Y => sample_out_0_sqmuxa);
    
    sample_out_val_RNO : NOR2A
      port map(A => sample_f1_val_0, B => un2_sample_in_val, Y
         => sample_out_val_4);
    
    \sample_out[53]\ : DFN1E1
      port map(D => sample_f1(85), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(42));
    
    \sample_out[28]\ : DFN1E1
      port map(D => sample_f1_wdata_67, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(67));
    
    \counter_RNO[27]\ : NOR2B
      port map(A => I_196_2, B => un2_sample_in_val, Y => 
        \counter_4[27]\);
    
    \sample_out[59]\ : DFN1E1
      port map(D => sample_f1(91), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(36));
    
    \counter_RNI0MBF1_1[10]\ : NOR3B
      port map(A => sample_f1_val_0, B => HRESETn_c, C => 
        un2_sample_in_val_0, Y => sample_out_0_sqmuxa_2);
    
    un3_counter_I_192 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[22]\, Y => \DWACT_FDEC_E[23]\);
    
    \sample_out[24]\ : DFN1E1
      port map(D => sample_f1_wdata_71, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(71));
    
    un3_counter_I_55 : OR3
      port map(A => \DWACT_FDEC_E[4]\, B => \counter[8]_net_1\, C
         => \counter[9]_net_1\, Y => N_103);
    
    \sample_out[42]\ : DFN1E1
      port map(D => sample_f1_wdata_53, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(53));
    
    un3_counter_I_118 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[13]\);
    
    \sample_out[40]\ : DFN1E1
      port map(D => sample_f1_wdata_55, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(55));
    
    \sample_out[83]\ : DFN1E1
      port map(D => sample_f1_wdata_12, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(12));
    
    \sample_out[89]\ : DFN1E1
      port map(D => sample_f1_wdata_6, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(6));
    
    \counter_RNIV507[8]\ : NOR2
      port map(A => \counter[8]_net_1\, B => \counter[9]_net_1\, 
        Y => un2_sample_in_val_9);
    
    un3_counter_I_189 : OR3
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        C => \counter[26]_net_1\, Y => \DWACT_FDEC_E[22]\);
    
    \counter_RNO[24]\ : NOR2B
      port map(A => I_166_2, B => un2_sample_in_val, Y => 
        \counter_4[24]\);
    
    \counter[7]\ : DFN1E1C0
      port map(D => I_38_2, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f1_val, Q => \counter[7]_net_1\);
    
    un3_counter_I_105 : XNOR2
      port map(A => N_68, B => \counter[17]_net_1\, Y => I_105_2);
    
    \sample_out[6]\ : DFN1E1
      port map(D => sample_f1_wdata_89, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(89));
    
    un3_counter_I_155 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[33]\, Y => N_32);
    
    un3_counter_I_179 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[20]\, Y => \DWACT_FDEC_E[21]\);
    
    \sample_out[62]\ : DFN1E1
      port map(D => sample_f1(94), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(33));
    
    \sample_out[60]\ : DFN1E1
      port map(D => sample_f1(92), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(35));
    
    un3_counter_I_65 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \counter[9]_net_1\, C
         => \counter[10]_net_1\, Y => N_96);
    
    \sample_out[35]\ : DFN1E1
      port map(D => sample_f1_wdata_60, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(60));
    
    \sample_out[91]\ : DFN1E1
      port map(D => sample_f1_wdata_4, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(4));
    
    un3_counter_I_135 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[15]\, Y => N_46);
    
    un3_counter_I_80 : OR2
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        Y => \DWACT_FDEC_E[8]\);
    
    \counter_RNIAEQF[20]\ : NOR3C
      port map(A => un2_sample_in_val_15, B => 
        un2_sample_in_val_14, C => un2_sample_in_val_20, Y => 
        un2_sample_in_val_24);
    
    un3_counter_I_16 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[0]\);
    
    \counter_RNO[20]\ : NOR2B
      port map(A => I_129_2, B => un2_sample_in_val, Y => 
        \counter_4[20]\);
    
    \sample_out[37]\ : DFN1E1
      port map(D => sample_f1_wdata_58, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(58));
    
    \sample_out[23]\ : DFN1E1
      port map(D => sample_f1_wdata_72, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(72));
    
    \sample_out[52]\ : DFN1E1
      port map(D => sample_f1(84), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(43));
    
    \sample_out[29]\ : DFN1E1
      port map(D => sample_f1_wdata_66, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(66));
    
    \counter_RNI3C64[22]\ : NOR3A
      port map(A => un2_sample_in_val_7, B => \counter[22]_net_1\, 
        C => \counter[19]_net_1\, Y => un2_sample_in_val_17);
    
    un3_counter_I_76 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \counter[12]_net_1\, Y => N_88);
    
    un3_counter_I_30 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[1]\, C
         => \counter[5]_net_1\, Y => N_121);
    
    \sample_out[50]\ : DFN1E1
      port map(D => sample_f1(82), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(45));
    
    \sample_out[18]\ : DFN1E1
      port map(D => sample_f1_wdata_77, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(77));
    
    \sample_out[9]\ : DFN1E1
      port map(D => sample_f1_wdata_86, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(86));
    
    \sample_out[7]\ : DFN1E1
      port map(D => sample_f1_wdata_88, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(88));
    
    \sample_out[78]\ : DFN1E1
      port map(D => sample_f1(110), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(17));
    
    un3_counter_I_83 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[8]\, Y => N_83);
    
    un3_counter_I_19 : OR2
      port map(A => \counter[3]_net_1\, B => \DWACT_FDEC_E[0]\, Y
         => N_129);
    
    \sample_out[14]\ : DFN1E1
      port map(D => sample_f1_wdata_81, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f3_wdata(81));
    
    \sample_out[82]\ : DFN1E1
      port map(D => sample_f1_wdata_13, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(13));
    
    \counter[9]\ : DFN1E1C0
      port map(D => \counter_4[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[9]_net_1\);
    
    \sample_out[74]\ : DFN1E1
      port map(D => sample_f1(106), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f3_wdata(21));
    
    \sample_out[80]\ : DFN1E1
      port map(D => sample_f1_wdata_15, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(15));
    
    \counter_RNIKN371_0[10]\ : OR3C
      port map(A => un2_sample_in_val_23, B => 
        un2_sample_in_val_22, C => un2_sample_in_val_24, Y => 
        un2_sample_in_val);
    
    \counter_RNO[19]\ : NOR2B
      port map(A => I_122_2, B => un2_sample_in_val, Y => 
        \counter_4[19]\);
    
    un3_counter_I_152 : OR3
      port map(A => \DWACT_FDEC_E[34]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[29]\);
    
    \counter_RNO[9]\ : NOR2B
      port map(A => I_52_2, B => un2_sample_in_val_0, Y => 
        \counter_4[9]\);
    
    \counter_RNIQKE[21]\ : NOR2
      port map(A => \counter[18]_net_1\, B => \counter[21]_net_1\, 
        Y => un2_sample_in_val_11);
    
    \counter[8]\ : DFN1E1C0
      port map(D => \counter_4[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[8]_net_1\);
    
    un3_counter_I_84 : XNOR2
      port map(A => N_83, B => \counter[14]_net_1\, Y => I_84_2);
    
    un3_counter_I_143 : XNOR2
      port map(A => N_41, B => \counter[22]_net_1\, Y => I_143_2);
    
    \counter[18]\ : DFN1E1C0
      port map(D => \counter_4[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f1_val, Q => \counter[18]_net_1\);
    
    un3_counter_I_90 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[9]\, Y => N_78);
    
    un3_counter_I_169 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \counter[24]_net_1\, Y => \DWACT_FDEC_E[19]\);
    
    un3_counter_I_132 : OR3
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        C => \counter[20]_net_1\, Y => \DWACT_FDEC_E[15]\);
    
    \sample_out[8]\ : DFN1E1
      port map(D => sample_f1_wdata_87, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f3_wdata(87));
    
    \sample_out[41]\ : DFN1E1
      port map(D => sample_f1_wdata_54, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(54));
    
    \counter_RNO[16]\ : NOR2B
      port map(A => I_98_2, B => un2_sample_in_val_0, Y => 
        \counter_4[16]\);
    
    \counter[0]\ : DFN1E1C0
      port map(D => I_4_2, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f1_val_0, Q => \counter[0]_net_1\);
    
    \sample_out[46]\ : DFN1E1
      port map(D => sample_f1_wdata_49, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(49));
    
    \counter_RNIKDT[27]\ : NOR3A
      port map(A => un2_sample_in_val_1, B => \counter[11]_net_1\, 
        C => \counter[27]_net_1\, Y => un2_sample_in_val_14);
    
    \sample_out[3]\ : DFN1E1
      port map(D => sample_f1_wdata_92, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1, Q => sample_f3_wdata(92));
    
    un3_counter_I_34 : OR3
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        C => \counter[5]_net_1\, Y => \DWACT_FDEC_E[2]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Downsampling_6_16_96 is

    port( sample_f0             : in    std_logic_vector(111 downto 80);
          sample_f0_wdata_95    : in    std_logic;
          sample_f0_wdata_94    : in    std_logic;
          sample_f0_wdata_93    : in    std_logic;
          sample_f0_wdata_92    : in    std_logic;
          sample_f0_wdata_91    : in    std_logic;
          sample_f0_wdata_90    : in    std_logic;
          sample_f0_wdata_89    : in    std_logic;
          sample_f0_wdata_88    : in    std_logic;
          sample_f0_wdata_87    : in    std_logic;
          sample_f0_wdata_86    : in    std_logic;
          sample_f0_wdata_85    : in    std_logic;
          sample_f0_wdata_84    : in    std_logic;
          sample_f0_wdata_83    : in    std_logic;
          sample_f0_wdata_82    : in    std_logic;
          sample_f0_wdata_81    : in    std_logic;
          sample_f0_wdata_80    : in    std_logic;
          sample_f0_wdata_79    : in    std_logic;
          sample_f0_wdata_78    : in    std_logic;
          sample_f0_wdata_77    : in    std_logic;
          sample_f0_wdata_76    : in    std_logic;
          sample_f0_wdata_75    : in    std_logic;
          sample_f0_wdata_74    : in    std_logic;
          sample_f0_wdata_73    : in    std_logic;
          sample_f0_wdata_72    : in    std_logic;
          sample_f0_wdata_71    : in    std_logic;
          sample_f0_wdata_70    : in    std_logic;
          sample_f0_wdata_69    : in    std_logic;
          sample_f0_wdata_68    : in    std_logic;
          sample_f0_wdata_67    : in    std_logic;
          sample_f0_wdata_66    : in    std_logic;
          sample_f0_wdata_65    : in    std_logic;
          sample_f0_wdata_64    : in    std_logic;
          sample_f0_wdata_63    : in    std_logic;
          sample_f0_wdata_62    : in    std_logic;
          sample_f0_wdata_61    : in    std_logic;
          sample_f0_wdata_60    : in    std_logic;
          sample_f0_wdata_59    : in    std_logic;
          sample_f0_wdata_58    : in    std_logic;
          sample_f0_wdata_57    : in    std_logic;
          sample_f0_wdata_56    : in    std_logic;
          sample_f0_wdata_55    : in    std_logic;
          sample_f0_wdata_54    : in    std_logic;
          sample_f0_wdata_53    : in    std_logic;
          sample_f0_wdata_52    : in    std_logic;
          sample_f0_wdata_51    : in    std_logic;
          sample_f0_wdata_50    : in    std_logic;
          sample_f0_wdata_49    : in    std_logic;
          sample_f0_wdata_48    : in    std_logic;
          sample_f0_wdata_15    : in    std_logic;
          sample_f0_wdata_14    : in    std_logic;
          sample_f0_wdata_13    : in    std_logic;
          sample_f0_wdata_12    : in    std_logic;
          sample_f0_wdata_11    : in    std_logic;
          sample_f0_wdata_10    : in    std_logic;
          sample_f0_wdata_9     : in    std_logic;
          sample_f0_wdata_8     : in    std_logic;
          sample_f0_wdata_7     : in    std_logic;
          sample_f0_wdata_6     : in    std_logic;
          sample_f0_wdata_5     : in    std_logic;
          sample_f0_wdata_4     : in    std_logic;
          sample_f0_wdata_3     : in    std_logic;
          sample_f0_wdata_2     : in    std_logic;
          sample_f0_wdata_1     : in    std_logic;
          sample_f0_wdata_0     : in    std_logic;
          sample_f2_wdata       : out   std_logic_vector(95 downto 0);
          sample_f0_val         : in    std_logic;
          sample_f0_val_1       : in    std_logic;
          HRESETn_c             : in    std_logic;
          HCLK_c                : in    std_logic;
          sample_f2_val         : out   std_logic;
          sample_f0_val_0       : in    std_logic;
          sample_out_0_sqmuxa_1 : in    std_logic
        );

end Downsampling_6_16_96;

architecture DEF_ARCH of Downsampling_6_16_96 is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal un6_sample_in_val_24_0, un6_sample_in_val_15, 
        un6_sample_in_val_14, un6_sample_in_val_20, 
        un6_sample_in_val_25_0, un6_sample_in_val_17, 
        un6_sample_in_val_16, un6_sample_in_val_23, 
        sample_out_0_sqmuxa_2, sample_out_0_sqmuxa_1_0, 
        sample_out_0_sqmuxa_0, N_137, \counter[1]_net_1\, 
        \counter[0]_net_1\, N_129, \counter[3]_net_1\, 
        \DWACT_FDEC_E[0]\, N_106, \counter[8]_net_1\, 
        \DWACT_FDEC_E[4]\, N_91, \DWACT_FDEC_E[7]\, 
        \DWACT_FDEC_E[6]\, un6_sample_in_val_25, 
        un6_sample_in_val_24, un6_sample_in_val_9, 
        un6_sample_in_val_8, un6_sample_in_val_19, 
        un6_sample_in_val_13, \counter[24]_net_1\, 
        un6_sample_in_val_11, \counter[15]_net_1\, 
        \counter[12]_net_1\, un6_sample_in_val_7, 
        \counter[22]_net_1\, \counter[19]_net_1\, 
        un6_sample_in_val_5, \counter[10]_net_1\, 
        \counter[7]_net_1\, un6_sample_in_val_3, 
        \counter[23]_net_1\, \counter[20]_net_1\, 
        un6_sample_in_val_1, \counter[11]_net_1\, 
        \counter[27]_net_1\, \counter[18]_net_1\, 
        \counter[21]_net_1\, \counter[9]_net_1\, 
        \counter[4]_net_1\, \counter[6]_net_1\, 
        \counter[25]_net_1\, \counter[2]_net_1\, 
        \counter[13]_net_1\, \counter[16]_net_1\, 
        \counter[26]_net_1\, \counter[5]_net_1\, 
        \counter[14]_net_1\, \counter[17]_net_1\, 
        sample_out_val_9, \counter_4[5]\, I_24_1, \counter_4[7]\, 
        I_38_1, \counter_4[8]\, I_45_1, \counter_4[9]\, I_52_1, 
        \counter_4[10]\, I_56_1, \counter_4[11]\, I_66_1, 
        \counter_4[12]\, I_73_1, \counter_4[13]\, I_77_1, 
        \counter_4[14]\, I_84_1, \counter_4[15]\, I_91_1, 
        \counter_4[16]\, I_98_1, \counter_4[17]\, I_105_1, 
        \counter_4[18]\, I_115_1, \counter_4[19]\, I_122_1, 
        \counter_4[20]\, I_129_1, \counter_4[21]\, I_136_1, 
        \counter_4[22]\, I_143_1, \counter_4[23]\, I_156_1, 
        \counter_4[24]\, I_166_1, \counter_4[25]\, I_173_1, 
        \counter_4[26]\, I_186_1, \counter_4[27]\, I_196_1, 
        sample_out_0_sqmuxa, I_4_1, I_5_1, I_9_1, I_13_1, I_20_1, 
        I_31_2, N_4, \DWACT_FDEC_E[29]\, \DWACT_FDEC_E[30]\, 
        \DWACT_FDEC_E[23]\, \DWACT_FDEC_E[15]\, 
        \DWACT_FDEC_E[17]\, \DWACT_FDEC_E[22]\, N_11, 
        \DWACT_FDEC_E[21]\, \DWACT_FDEC_E[9]\, \DWACT_FDEC_E[12]\, 
        \DWACT_FDEC_E[20]\, N_20, \DWACT_FDEC_E[13]\, 
        \DWACT_FDEC_E[19]\, N_25, \DWACT_FDEC_E[18]\, N_32, 
        \DWACT_FDEC_E[33]\, \DWACT_FDEC_E[34]\, \DWACT_FDEC_E[2]\, 
        \DWACT_FDEC_E[5]\, N_41, \DWACT_FDEC_E[28]\, 
        \DWACT_FDEC_E[16]\, N_46, N_51, \DWACT_FDEC_E[14]\, N_56, 
        N_61, \DWACT_FDEC_E[10]\, N_68, \DWACT_FDEC_E[11]\, N_73, 
        N_78, N_83, \DWACT_FDEC_E[8]\, N_88, N_96, N_103, 
        \DWACT_FDEC_E[3]\, N_111, N_116, N_121, \DWACT_FDEC_E[1]\, 
        N_126, N_134, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \counter[19]\ : DFN1E1C0
      port map(D => \counter_4[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[19]_net_1\);
    
    \sample_out[22]\ : DFN1E1
      port map(D => sample_f0_wdata_73, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(73));
    
    \sample_out[20]\ : DFN1E1
      port map(D => sample_f0_wdata_75, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(75));
    
    \sample_out[13]\ : DFN1E1
      port map(D => sample_f0_wdata_82, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(82));
    
    \sample_out[1]\ : DFN1E1
      port map(D => sample_f0_wdata_94, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(94));
    
    \sample_out[19]\ : DFN1E1
      port map(D => sample_f0_wdata_76, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(76));
    
    un3_counter_I_142 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[16]\, Y => N_41);
    
    \sample_out[61]\ : DFN1E1
      port map(D => sample_f0(93), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(34));
    
    \sample_out[66]\ : DFN1E1
      port map(D => sample_f0(98), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(29));
    
    \sample_out[73]\ : DFN1E1
      port map(D => sample_f0(105), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(22));
    
    \sample_out[79]\ : DFN1E1
      port map(D => sample_f0(111), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(16));
    
    \sample_out[38]\ : DFN1E1
      port map(D => sample_f0_wdata_57, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(57));
    
    un3_counter_I_27 : OR2
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        Y => \DWACT_FDEC_E[1]\);
    
    \sample_out[95]\ : DFN1E1
      port map(D => sample_f0_wdata_0, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(0));
    
    \counter_RNO[11]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_66_1, Y => \counter_4[11]\);
    
    \counter_RNISF54[20]\ : NOR3A
      port map(A => un6_sample_in_val_3, B => \counter[23]_net_1\, 
        C => \counter[20]_net_1\, Y => un6_sample_in_val_15);
    
    \counter_RNID1T[12]\ : NOR3A
      port map(A => un6_sample_in_val_11, B => 
        \counter[15]_net_1\, C => \counter[12]_net_1\, Y => 
        un6_sample_in_val_19);
    
    \sample_out[34]\ : DFN1E1
      port map(D => sample_f0_wdata_61, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(61));
    
    un3_counter_I_4 : INV
      port map(A => \counter[0]_net_1\, Y => I_4_1);
    
    \counter[11]\ : DFN1E1C0
      port map(D => \counter_4[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[11]_net_1\);
    
    un3_counter_I_94 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, Y
         => \DWACT_FDEC_E[10]\);
    
    un3_counter_I_186 : XNOR2
      port map(A => N_11, B => \counter[26]_net_1\, Y => I_186_1);
    
    \counter_RNO[15]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_91_1, Y => \counter_4[15]\);
    
    un3_counter_I_108 : OR3
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        C => \counter[17]_net_1\, Y => \DWACT_FDEC_E[12]\);
    
    un3_counter_I_121 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \counter[18]_net_1\, Y => N_56);
    
    \sample_out[51]\ : DFN1E1
      port map(D => sample_f0(83), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(44));
    
    \sample_out[56]\ : DFN1E1
      port map(D => sample_f0(88), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(39));
    
    un3_counter_I_176 : OR2
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        Y => \DWACT_FDEC_E[20]\);
    
    \sample_out[0]\ : DFN1E1
      port map(D => sample_f0_wdata_95, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(95));
    
    \counter_RNO[7]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_38_1, Y => \counter_4[7]\);
    
    \counter[6]\ : DFN1E1C0
      port map(D => I_31_2, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f0_val, Q => \counter[6]_net_1\);
    
    un3_counter_I_48 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => \DWACT_FDEC_E[4]\);
    
    un3_counter_I_114 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[10]\, 
        C => \DWACT_FDEC_E[12]\, Y => N_61);
    
    \counter_RNIPSE[14]\ : NOR2
      port map(A => \counter[14]_net_1\, B => \counter[17]_net_1\, 
        Y => un6_sample_in_val_1);
    
    \counter[21]\ : DFN1E1C0
      port map(D => \counter_4[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[21]_net_1\);
    
    un3_counter_I_13 : XNOR2
      port map(A => N_134, B => \counter[3]_net_1\, Y => I_13_1);
    
    \counter_RNIF507[3]\ : NOR2
      port map(A => \counter[3]_net_1\, B => \counter[0]_net_1\, 
        Y => un6_sample_in_val_13);
    
    \counter_RNI3LBF1_1[10]\ : NOR3C
      port map(A => un6_sample_in_val_24_0, B => 
        un6_sample_in_val_25_0, C => sample_out_0_sqmuxa_1, Y => 
        sample_out_0_sqmuxa_2);
    
    \sample_out[81]\ : DFN1E1
      port map(D => sample_f0_wdata_14, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(14));
    
    \sample_out[86]\ : DFN1E1
      port map(D => sample_f0_wdata_9, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(9));
    
    \counter_RNIOKE[21]\ : NOR2
      port map(A => \counter[18]_net_1\, B => \counter[21]_net_1\, 
        Y => un6_sample_in_val_11);
    
    \counter[3]\ : DFN1E1C0
      port map(D => I_13_1, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f0_val, Q => \counter[3]_net_1\);
    
    \counter[2]\ : DFN1E1C0
      port map(D => I_9_1, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f0_val, Q => \counter[2]_net_1\);
    
    un3_counter_I_73 : XNOR2
      port map(A => N_91, B => \counter[12]_net_1\, Y => I_73_1);
    
    \counter_RNO[8]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_45_1, Y => \counter_4[8]\);
    
    \counter_RNIUDQF[20]\ : NOR3C
      port map(A => un6_sample_in_val_15, B => 
        un6_sample_in_val_14, C => un6_sample_in_val_20, Y => 
        un6_sample_in_val_24_0);
    
    \counter_RNO[13]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_77_1, Y => \counter_4[13]\);
    
    un3_counter_I_52 : XNOR2
      port map(A => N_106, B => \counter[9]_net_1\, Y => I_52_1);
    
    \sample_out[12]\ : DFN1E1
      port map(D => sample_f0_wdata_83, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(83));
    
    \counter_RNIQ89N[10]\ : NOR3C
      port map(A => un6_sample_in_val_17, B => 
        un6_sample_in_val_16, C => un6_sample_in_val_23, Y => 
        un6_sample_in_val_25_0);
    
    \sample_out[10]\ : DFN1E1
      port map(D => sample_f0_wdata_85, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(85));
    
    \sample_out[45]\ : DFN1E1
      port map(D => sample_f0_wdata_50, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(50));
    
    \counter_RNO[12]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_73_1, Y => \counter_4[12]\);
    
    \counter_RNIT507[8]\ : NOR2
      port map(A => \counter[8]_net_1\, B => \counter[9]_net_1\, 
        Y => un6_sample_in_val_9);
    
    \sample_out[72]\ : DFN1E1
      port map(D => sample_f0(104), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(23));
    
    \sample_out[33]\ : DFN1E1
      port map(D => sample_f0_wdata_62, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(62));
    
    \sample_out[39]\ : DFN1E1
      port map(D => sample_f0_wdata_56, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(56));
    
    \counter[17]\ : DFN1E1C0
      port map(D => \counter_4[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[17]_net_1\);
    
    \sample_out[70]\ : DFN1E1
      port map(D => sample_f0(102), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(25));
    
    un3_counter_I_41 : OR2
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        Y => \DWACT_FDEC_E[3]\);
    
    un3_counter_I_159 : OR3
      port map(A => \counter[21]_net_1\, B => \counter[22]_net_1\, 
        C => \counter[23]_net_1\, Y => \DWACT_FDEC_E[17]\);
    
    \counter[4]\ : DFN1E1C0
      port map(D => I_20_1, CLK => HCLK_c, CLR => HRESETn_c, E
         => sample_f0_val, Q => \counter[4]_net_1\);
    
    un3_counter_I_5 : XNOR2
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        Y => I_5_1);
    
    \counter_RNIGDT[27]\ : NOR3A
      port map(A => un6_sample_in_val_1, B => \counter[11]_net_1\, 
        C => \counter[27]_net_1\, Y => un6_sample_in_val_14);
    
    un3_counter_I_125 : OR2
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        Y => \DWACT_FDEC_E[14]\);
    
    \counter[10]\ : DFN1E1C0
      port map(D => \counter_4[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[10]_net_1\);
    
    \sample_out[5]\ : DFN1E1
      port map(D => sample_f0_wdata_90, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(90));
    
    \sample_out[47]\ : DFN1E1
      port map(D => sample_f0_wdata_48, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(48));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter[13]\ : DFN1E1C0
      port map(D => \counter_4[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[13]_net_1\);
    
    un3_counter_I_62 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[6]\);
    
    \sample_out[65]\ : DFN1E1
      port map(D => sample_f0(97), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(30));
    
    un3_counter_I_139 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        Y => \DWACT_FDEC_E[16]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sample_out[21]\ : DFN1E1
      port map(D => sample_f0_wdata_74, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(74));
    
    \counter[12]\ : DFN1E1C0
      port map(D => \counter_4[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[12]_net_1\);
    
    \sample_out[26]\ : DFN1E1
      port map(D => sample_f0_wdata_69, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(69));
    
    \sample_out[2]\ : DFN1E1
      port map(D => sample_f0_wdata_93, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(93));
    
    \counter[27]\ : DFN1E1C0
      port map(D => \counter_4[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[27]_net_1\);
    
    un3_counter_I_111 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[28]\);
    
    \sample_out[67]\ : DFN1E1
      port map(D => sample_f0(99), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(28));
    
    \counter[20]\ : DFN1E1C0
      port map(D => \counter_4[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[20]_net_1\);
    
    \sample_out[94]\ : DFN1E1
      port map(D => sample_f0_wdata_1, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(1));
    
    un3_counter_I_166 : XNOR2
      port map(A => N_25, B => \counter[24]_net_1\, Y => I_166_1);
    
    \counter_RNO[17]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_105_1, Y => \counter_4[17]\);
    
    \counter[23]\ : DFN1E1C0
      port map(D => \counter_4[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[23]_net_1\);
    
    un3_counter_I_149 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[34]\);
    
    \sample_out[55]\ : DFN1E1
      port map(D => sample_f0(87), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(40));
    
    \counter[22]\ : DFN1E1C0
      port map(D => \counter_4[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[22]_net_1\);
    
    \counter[15]\ : DFN1E1C0
      port map(D => \counter_4[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[15]_net_1\);
    
    un3_counter_I_8 : OR2
      port map(A => \counter[1]_net_1\, B => \counter[0]_net_1\, 
        Y => N_137);
    
    un3_counter_I_185 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[21]\, Y => N_11);
    
    un3_counter_I_196 : XNOR2
      port map(A => N_4, B => \counter[27]_net_1\, Y => I_196_1);
    
    \sample_out[32]\ : DFN1E1
      port map(D => sample_f0_wdata_63, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(63));
    
    un3_counter_I_51 : OR2
      port map(A => \counter[8]_net_1\, B => \DWACT_FDEC_E[4]\, Y
         => N_106);
    
    un3_counter_I_122 : XNOR2
      port map(A => N_56, B => \counter[19]_net_1\, Y => I_122_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sample_out[57]\ : DFN1E1
      port map(D => sample_f0(89), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(38));
    
    \sample_out[30]\ : DFN1E1
      port map(D => sample_f0_wdata_65, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(65));
    
    \counter_RNO[14]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_84_1, Y => \counter_4[14]\);
    
    \sample_out[85]\ : DFN1E1
      port map(D => sample_f0_wdata_10, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(10));
    
    \counter[1]\ : DFN1E1C0
      port map(D => I_5_1, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f0_val, Q => \counter[1]_net_1\);
    
    \counter_RNO[26]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_186_1, Y => \counter_4[26]\);
    
    \sample_out[4]\ : DFN1E1
      port map(D => sample_f0_wdata_91, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(91));
    
    \counter_RNO[5]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_24_1, Y => \counter_4[5]\);
    
    \counter[25]\ : DFN1E1C0
      port map(D => \counter_4[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[25]_net_1\);
    
    sample_out_val : DFN1C0
      port map(D => sample_out_val_9, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f2_val);
    
    \sample_out[87]\ : DFN1E1
      port map(D => sample_f0_wdata_8, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(8));
    
    un3_counter_I_115 : XNOR2
      port map(A => N_61, B => \counter[18]_net_1\, Y => I_115_1);
    
    \counter_RNIUDQF_0[20]\ : NOR3C
      port map(A => un6_sample_in_val_15, B => 
        un6_sample_in_val_14, C => un6_sample_in_val_20, Y => 
        un6_sample_in_val_24);
    
    un3_counter_I_87 : OR3
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        C => \counter[14]_net_1\, Y => \DWACT_FDEC_E[9]\);
    
    un3_counter_I_173 : XNOR2
      port map(A => N_20, B => \counter[25]_net_1\, Y => I_173_1);
    
    \sample_out[48]\ : DFN1E1
      port map(D => sample_f0(80), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(47));
    
    un3_counter_I_38 : XNOR2
      port map(A => N_116, B => \counter[7]_net_1\, Y => I_38_1);
    
    \sample_out[93]\ : DFN1E1
      port map(D => sample_f0_wdata_2, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(2));
    
    \sample_out[11]\ : DFN1E1
      port map(D => sample_f0_wdata_84, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(84));
    
    \sample_out[16]\ : DFN1E1
      port map(D => sample_f0_wdata_79, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(79));
    
    \counter[5]\ : DFN1E1C0
      port map(D => \counter_4[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[5]_net_1\);
    
    \sample_out[44]\ : DFN1E1
      port map(D => sample_f0_wdata_51, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(51));
    
    \sample_out[71]\ : DFN1E1
      port map(D => sample_f0(103), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(24));
    
    \counter_RNI0DTE[12]\ : NOR3C
      port map(A => un6_sample_in_val_9, B => un6_sample_in_val_8, 
        C => un6_sample_in_val_19, Y => un6_sample_in_val_23);
    
    \sample_out[76]\ : DFN1E1
      port map(D => sample_f0(108), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(19));
    
    \counter_RNI3LBF1_0[10]\ : NOR3C
      port map(A => un6_sample_in_val_24_0, B => 
        un6_sample_in_val_25_0, C => sample_out_0_sqmuxa_1, Y => 
        sample_out_0_sqmuxa_0);
    
    un3_counter_I_37 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \counter[6]_net_1\, Y => N_116);
    
    \counter_RNO[10]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_56_1, Y => \counter_4[10]\);
    
    un3_counter_I_9 : XNOR2
      port map(A => N_137, B => \counter[2]_net_1\, Y => I_9_1);
    
    \counter_RNO[21]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_136_1, Y => \counter_4[21]\);
    
    un3_counter_I_20 : XNOR2
      port map(A => N_129, B => \counter[4]_net_1\, Y => I_20_1);
    
    un3_counter_I_182 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[30]\);
    
    \sample_out[68]\ : DFN1E1
      port map(D => sample_f0(100), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(27));
    
    \sample_out[25]\ : DFN1E1
      port map(D => sample_f0_wdata_70, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(70));
    
    un3_counter_I_56 : XNOR2
      port map(A => N_103, B => \counter[10]_net_1\, Y => I_56_1);
    
    \counter_RNIM507[4]\ : NOR2
      port map(A => \counter[4]_net_1\, B => \counter[6]_net_1\, 
        Y => un6_sample_in_val_8);
    
    \counter[16]\ : DFN1E1C0
      port map(D => \counter_4[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[16]_net_1\);
    
    \counter_RNO[25]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_173_1, Y => \counter_4[25]\);
    
    un3_counter_I_172 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[19]\, Y => N_20);
    
    un3_counter_I_104 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \DWACT_FDEC_E[11]\, Y => N_68);
    
    \sample_out[64]\ : DFN1E1
      port map(D => sample_f0(96), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(31));
    
    un3_counter_I_31 : XNOR2
      port map(A => N_121, B => \counter[6]_net_1\, Y => I_31_2);
    
    un3_counter_I_98 : XNOR2
      port map(A => N_73, B => \counter[16]_net_1\, Y => I_98_1);
    
    un3_counter_I_23 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \counter[3]_net_1\, C
         => \counter[4]_net_1\, Y => N_126);
    
    \sample_out[27]\ : DFN1E1
      port map(D => sample_f0_wdata_68, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(68));
    
    un3_counter_I_59 : OR3
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        C => \counter[8]_net_1\, Y => \DWACT_FDEC_E[5]\);
    
    un3_counter_I_12 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => N_134);
    
    \counter_RNI3LBF1_2[10]\ : NOR3C
      port map(A => un6_sample_in_val_24_0, B => 
        un6_sample_in_val_25_0, C => sample_out_0_sqmuxa_1, Y => 
        sample_out_0_sqmuxa_1_0);
    
    un3_counter_I_165 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[18]\, Y => N_25);
    
    un3_counter_I_156 : XNOR2
      port map(A => N_32, B => \counter[23]_net_1\, Y => I_156_1);
    
    un3_counter_I_97 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \counter[15]_net_1\, Y => N_73);
    
    un3_counter_I_128 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[14]\, Y => N_51);
    
    \counter_RNIRF54[10]\ : NOR3A
      port map(A => un6_sample_in_val_5, B => \counter[10]_net_1\, 
        C => \counter[7]_net_1\, Y => un6_sample_in_val_16);
    
    un3_counter_I_72 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[6]\, Y
         => N_91);
    
    \sample_out[58]\ : DFN1E1
      port map(D => sample_f0(90), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(37));
    
    \counter[26]\ : DFN1E1C0
      port map(D => \counter_4[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[26]_net_1\);
    
    un3_counter_I_66 : XNOR2
      port map(A => N_96, B => \counter[11]_net_1\, Y => I_66_1);
    
    \counter_RNO[23]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_156_1, Y => \counter_4[23]\);
    
    \sample_out[54]\ : DFN1E1
      port map(D => sample_f0(86), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(41));
    
    \sample_out[43]\ : DFN1E1
      port map(D => sample_f0_wdata_52, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(52));
    
    \sample_out[49]\ : DFN1E1
      port map(D => sample_f0(81), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(46));
    
    \counter_RNI3LBF1[10]\ : NOR3C
      port map(A => un6_sample_in_val_24, B => 
        un6_sample_in_val_25, C => sample_out_0_sqmuxa_1, Y => 
        sample_out_0_sqmuxa);
    
    un3_counter_I_45 : XNOR2
      port map(A => N_111, B => \counter[8]_net_1\, Y => I_45_1);
    
    un3_counter_I_24 : XNOR2
      port map(A => N_126, B => \counter[5]_net_1\, Y => I_24_1);
    
    un3_counter_I_195 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[23]\, Y => N_4);
    
    \sample_out[92]\ : DFN1E1
      port map(D => sample_f0_wdata_3, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(3));
    
    \counter[14]\ : DFN1E1C0
      port map(D => \counter_4[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[14]_net_1\);
    
    un3_counter_I_136 : XNOR2
      port map(A => N_46, B => \counter[21]_net_1\, Y => I_136_1);
    
    \sample_out[88]\ : DFN1E1
      port map(D => sample_f0_wdata_7, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(7));
    
    \counter_RNIVB64[22]\ : NOR3A
      port map(A => un6_sample_in_val_7, B => \counter[22]_net_1\, 
        C => \counter[19]_net_1\, Y => un6_sample_in_val_17);
    
    \sample_out[90]\ : DFN1E1
      port map(D => sample_f0_wdata_5, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(5));
    
    un3_counter_I_91 : XNOR2
      port map(A => N_78, B => \counter[15]_net_1\, Y => I_91_1);
    
    \counter_RNO[22]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_143_1, Y => \counter_4[22]\);
    
    \sample_out[31]\ : DFN1E1
      port map(D => sample_f0_wdata_64, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(64));
    
    \sample_out[36]\ : DFN1E1
      port map(D => sample_f0_wdata_59, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(59));
    
    un3_counter_I_69 : OR3
      port map(A => \counter[9]_net_1\, B => \counter[10]_net_1\, 
        C => \counter[11]_net_1\, Y => \DWACT_FDEC_E[7]\);
    
    \sample_out[84]\ : DFN1E1
      port map(D => sample_f0_wdata_11, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(11));
    
    \sample_out[63]\ : DFN1E1
      port map(D => sample_f0(95), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(32));
    
    \sample_out[69]\ : DFN1E1
      port map(D => sample_f0(101), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(26));
    
    \sample_out[15]\ : DFN1E1
      port map(D => sample_f0_wdata_80, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(80));
    
    un3_counter_I_129 : XNOR2
      port map(A => N_51, B => \counter[20]_net_1\, Y => I_129_1);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un3_counter_I_146 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        C => \counter[22]_net_1\, Y => \DWACT_FDEC_E[33]\);
    
    \counter[24]\ : DFN1E1C0
      port map(D => \counter_4[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[24]_net_1\);
    
    un3_counter_I_101 : OR2
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        Y => \DWACT_FDEC_E[11]\);
    
    \sample_out[75]\ : DFN1E1
      port map(D => sample_f0(107), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(20));
    
    \counter_RNIIGNA[24]\ : NOR3A
      port map(A => un6_sample_in_val_13, B => \counter[1]_net_1\, 
        C => \counter[24]_net_1\, Y => un6_sample_in_val_20);
    
    \counter_RNI9JN3[26]\ : NOR2
      port map(A => \counter[26]_net_1\, B => \counter[5]_net_1\, 
        Y => un6_sample_in_val_3);
    
    un3_counter_I_162 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        Y => \DWACT_FDEC_E[18]\);
    
    \counter_RNIQ89N_0[10]\ : NOR3C
      port map(A => un6_sample_in_val_17, B => 
        un6_sample_in_val_16, C => un6_sample_in_val_23, Y => 
        un6_sample_in_val_25);
    
    un3_counter_I_77 : XNOR2
      port map(A => N_88, B => \counter[13]_net_1\, Y => I_77_1);
    
    \sample_out[17]\ : DFN1E1
      port map(D => sample_f0_wdata_78, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(78));
    
    \counter_RNO[18]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_115_1, Y => \counter_4[18]\);
    
    un3_counter_I_44 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => N_111);
    
    \sample_out[77]\ : DFN1E1
      port map(D => sample_f0(109), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(18));
    
    sample_out_val_RNO : NOR3C
      port map(A => un6_sample_in_val_24_0, B => 
        un6_sample_in_val_25_0, C => sample_f0_val_0, Y => 
        sample_out_val_9);
    
    \sample_out[53]\ : DFN1E1
      port map(D => sample_f0(85), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(42));
    
    \sample_out[28]\ : DFN1E1
      port map(D => sample_f0_wdata_67, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(67));
    
    \counter_RNO[27]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_196_1, Y => \counter_4[27]\);
    
    \sample_out[59]\ : DFN1E1
      port map(D => sample_f0(91), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(36));
    
    un3_counter_I_192 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[22]\, Y => \DWACT_FDEC_E[23]\);
    
    \sample_out[24]\ : DFN1E1
      port map(D => sample_f0_wdata_71, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(71));
    
    un3_counter_I_55 : OR3
      port map(A => \DWACT_FDEC_E[4]\, B => \counter[8]_net_1\, C
         => \counter[9]_net_1\, Y => N_103);
    
    \sample_out[42]\ : DFN1E1
      port map(D => sample_f0_wdata_53, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(53));
    
    un3_counter_I_118 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[13]\);
    
    \sample_out[40]\ : DFN1E1
      port map(D => sample_f0_wdata_55, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(55));
    
    \sample_out[83]\ : DFN1E1
      port map(D => sample_f0_wdata_12, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(12));
    
    \sample_out[89]\ : DFN1E1
      port map(D => sample_f0_wdata_6, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(6));
    
    un3_counter_I_189 : OR3
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        C => \counter[26]_net_1\, Y => \DWACT_FDEC_E[22]\);
    
    \counter_RNO[24]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_166_1, Y => \counter_4[24]\);
    
    \counter[7]\ : DFN1E1C0
      port map(D => \counter_4[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[7]_net_1\);
    
    un3_counter_I_105 : XNOR2
      port map(A => N_68, B => \counter[17]_net_1\, Y => I_105_1);
    
    \sample_out[6]\ : DFN1E1
      port map(D => sample_f0_wdata_89, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(89));
    
    un3_counter_I_155 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[33]\, Y => N_32);
    
    un3_counter_I_179 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[20]\, Y => \DWACT_FDEC_E[21]\);
    
    \sample_out[62]\ : DFN1E1
      port map(D => sample_f0(94), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(33));
    
    \counter_RNINKE[13]\ : NOR2
      port map(A => \counter[13]_net_1\, B => \counter[16]_net_1\, 
        Y => un6_sample_in_val_5);
    
    \sample_out[60]\ : DFN1E1
      port map(D => sample_f0(92), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(35));
    
    un3_counter_I_65 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \counter[9]_net_1\, C
         => \counter[10]_net_1\, Y => N_96);
    
    \sample_out[35]\ : DFN1E1
      port map(D => sample_f0_wdata_60, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(60));
    
    \sample_out[91]\ : DFN1E1
      port map(D => sample_f0_wdata_4, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(4));
    
    un3_counter_I_135 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[15]\, Y => N_46);
    
    un3_counter_I_80 : OR2
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        Y => \DWACT_FDEC_E[8]\);
    
    un3_counter_I_16 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[0]\);
    
    \counter_RNO[20]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_129_1, Y => \counter_4[20]\);
    
    \sample_out[37]\ : DFN1E1
      port map(D => sample_f0_wdata_58, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(58));
    
    \sample_out[23]\ : DFN1E1
      port map(D => sample_f0_wdata_72, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(72));
    
    \sample_out[52]\ : DFN1E1
      port map(D => sample_f0(84), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(43));
    
    \sample_out[29]\ : DFN1E1
      port map(D => sample_f0_wdata_66, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(66));
    
    un3_counter_I_76 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \counter[12]_net_1\, Y => N_88);
    
    un3_counter_I_30 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[1]\, C
         => \counter[5]_net_1\, Y => N_121);
    
    \sample_out[50]\ : DFN1E1
      port map(D => sample_f0(82), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(45));
    
    \sample_out[18]\ : DFN1E1
      port map(D => sample_f0_wdata_77, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(77));
    
    \sample_out[9]\ : DFN1E1
      port map(D => sample_f0_wdata_86, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(86));
    
    \sample_out[7]\ : DFN1E1
      port map(D => sample_f0_wdata_88, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(88));
    
    \sample_out[78]\ : DFN1E1
      port map(D => sample_f0(110), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(17));
    
    un3_counter_I_83 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[8]\, Y => N_83);
    
    un3_counter_I_19 : OR2
      port map(A => \counter[3]_net_1\, B => \DWACT_FDEC_E[0]\, Y
         => N_129);
    
    \sample_out[14]\ : DFN1E1
      port map(D => sample_f0_wdata_81, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f2_wdata(81));
    
    \sample_out[82]\ : DFN1E1
      port map(D => sample_f0_wdata_13, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(13));
    
    \counter[9]\ : DFN1E1C0
      port map(D => \counter_4[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[9]_net_1\);
    
    \sample_out[74]\ : DFN1E1
      port map(D => sample_f0(106), CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f2_wdata(21));
    
    \sample_out[80]\ : DFN1E1
      port map(D => sample_f0_wdata_15, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(15));
    
    \counter_RNO[19]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_122_1, Y => \counter_4[19]\);
    
    un3_counter_I_152 : OR3
      port map(A => \DWACT_FDEC_E[34]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[29]\);
    
    \counter_RNO[9]\ : AOI1B
      port map(A => un6_sample_in_val_25_0, B => 
        un6_sample_in_val_24_0, C => I_52_1, Y => \counter_4[9]\);
    
    \counter_RNI5FN3[25]\ : NOR2
      port map(A => \counter[25]_net_1\, B => \counter[2]_net_1\, 
        Y => un6_sample_in_val_7);
    
    \counter[8]\ : DFN1E1C0
      port map(D => \counter_4[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[8]_net_1\);
    
    un3_counter_I_84 : XNOR2
      port map(A => N_83, B => \counter[14]_net_1\, Y => I_84_1);
    
    un3_counter_I_143 : XNOR2
      port map(A => N_41, B => \counter[22]_net_1\, Y => I_143_1);
    
    \counter[18]\ : DFN1E1C0
      port map(D => \counter_4[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val, Q => \counter[18]_net_1\);
    
    un3_counter_I_90 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[9]\, Y => N_78);
    
    un3_counter_I_169 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \counter[24]_net_1\, Y => \DWACT_FDEC_E[19]\);
    
    un3_counter_I_132 : OR3
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        C => \counter[20]_net_1\, Y => \DWACT_FDEC_E[15]\);
    
    \sample_out[8]\ : DFN1E1
      port map(D => sample_f0_wdata_87, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f2_wdata(87));
    
    \sample_out[41]\ : DFN1E1
      port map(D => sample_f0_wdata_54, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(54));
    
    \counter_RNO[16]\ : AOI1B
      port map(A => un6_sample_in_val_25, B => 
        un6_sample_in_val_24, C => I_98_1, Y => \counter_4[16]\);
    
    \counter[0]\ : DFN1E1C0
      port map(D => I_4_1, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f0_val_1, Q => \counter[0]_net_1\);
    
    \sample_out[46]\ : DFN1E1
      port map(D => sample_f0_wdata_49, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(49));
    
    \sample_out[3]\ : DFN1E1
      port map(D => sample_f0_wdata_92, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f2_wdata(92));
    
    un3_counter_I_34 : OR3
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        C => \counter[5]_net_1\, Y => \DWACT_FDEC_E[2]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1 is

    port( sample_f1_wdata_95 : in    std_logic;
          sample_f1_wdata_94 : in    std_logic;
          sample_f1_wdata_93 : in    std_logic;
          sample_f1_wdata_92 : in    std_logic;
          sample_f1_wdata_91 : in    std_logic;
          sample_f1_wdata_90 : in    std_logic;
          sample_f1_wdata_89 : in    std_logic;
          sample_f1_wdata_88 : in    std_logic;
          sample_f1_wdata_87 : in    std_logic;
          sample_f1_wdata_86 : in    std_logic;
          sample_f1_wdata_85 : in    std_logic;
          sample_f1_wdata_84 : in    std_logic;
          sample_f1_wdata_83 : in    std_logic;
          sample_f1_wdata_82 : in    std_logic;
          sample_f1_wdata_81 : in    std_logic;
          sample_f1_wdata_80 : in    std_logic;
          sample_f1_wdata_79 : in    std_logic;
          sample_f1_wdata_78 : in    std_logic;
          sample_f1_wdata_77 : in    std_logic;
          sample_f1_wdata_76 : in    std_logic;
          sample_f1_wdata_75 : in    std_logic;
          sample_f1_wdata_74 : in    std_logic;
          sample_f1_wdata_73 : in    std_logic;
          sample_f1_wdata_72 : in    std_logic;
          sample_f1_wdata_71 : in    std_logic;
          sample_f1_wdata_70 : in    std_logic;
          sample_f1_wdata_69 : in    std_logic;
          sample_f1_wdata_68 : in    std_logic;
          sample_f1_wdata_67 : in    std_logic;
          sample_f1_wdata_66 : in    std_logic;
          sample_f1_wdata_65 : in    std_logic;
          sample_f1_wdata_64 : in    std_logic;
          sample_f1_wdata_63 : in    std_logic;
          sample_f1_wdata_62 : in    std_logic;
          sample_f1_wdata_61 : in    std_logic;
          sample_f1_wdata_60 : in    std_logic;
          sample_f1_wdata_59 : in    std_logic;
          sample_f1_wdata_58 : in    std_logic;
          sample_f1_wdata_57 : in    std_logic;
          sample_f1_wdata_56 : in    std_logic;
          sample_f1_wdata_55 : in    std_logic;
          sample_f1_wdata_54 : in    std_logic;
          sample_f1_wdata_53 : in    std_logic;
          sample_f1_wdata_52 : in    std_logic;
          sample_f1_wdata_51 : in    std_logic;
          sample_f1_wdata_50 : in    std_logic;
          sample_f1_wdata_49 : in    std_logic;
          sample_f1_wdata_48 : in    std_logic;
          sample_f1_wdata_15 : in    std_logic;
          sample_f1_wdata_14 : in    std_logic;
          sample_f1_wdata_13 : in    std_logic;
          sample_f1_wdata_12 : in    std_logic;
          sample_f1_wdata_11 : in    std_logic;
          sample_f1_wdata_10 : in    std_logic;
          sample_f1_wdata_9  : in    std_logic;
          sample_f1_wdata_8  : in    std_logic;
          sample_f1_wdata_7  : in    std_logic;
          sample_f1_wdata_6  : in    std_logic;
          sample_f1_wdata_5  : in    std_logic;
          sample_f1_wdata_4  : in    std_logic;
          sample_f1_wdata_3  : in    std_logic;
          sample_f1_wdata_2  : in    std_logic;
          sample_f1_wdata_1  : in    std_logic;
          sample_f1_wdata_0  : in    std_logic;
          data_f1_out        : out   std_logic_vector(159 downto 64);
          nb_snapshot_param  : in    std_logic_vector(0 to 0);
          sample_f1_37       : in    std_logic;
          sample_f1_5        : in    std_logic;
          sample_f1_38       : in    std_logic;
          sample_f1_6        : in    std_logic;
          sample_f1_39       : in    std_logic;
          sample_f1_7        : in    std_logic;
          sample_f1_40       : in    std_logic;
          sample_f1_8        : in    std_logic;
          sample_f1_41       : in    std_logic;
          sample_f1_9        : in    std_logic;
          sample_f1_42       : in    std_logic;
          sample_f1_10       : in    std_logic;
          sample_f1_43       : in    std_logic;
          sample_f1_11       : in    std_logic;
          sample_f1_61       : in    std_logic;
          sample_f1_62       : in    std_logic;
          sample_f1_63       : in    std_logic;
          sample_f1_32       : in    std_logic;
          sample_f1_0        : in    std_logic;
          sample_f1_33       : in    std_logic;
          sample_f1_1        : in    std_logic;
          sample_f1_34       : in    std_logic;
          sample_f1_2        : in    std_logic;
          sample_f1_35       : in    std_logic;
          sample_f1_3        : in    std_logic;
          sample_f1_36       : in    std_logic;
          sample_f1_4        : in    std_logic;
          sample_f1_48       : in    std_logic;
          sample_f1_49       : in    std_logic;
          sample_f1_50       : in    std_logic;
          sample_f1_51       : in    std_logic;
          sample_f1_52       : in    std_logic;
          sample_f1_53       : in    std_logic;
          sample_f1_54       : in    std_logic;
          sample_f1_55       : in    std_logic;
          sample_f1_56       : in    std_logic;
          sample_f1_57       : in    std_logic;
          sample_f1_58       : in    std_logic;
          sample_f1_59       : in    std_logic;
          sample_f1_60       : in    std_logic;
          sample_f1_44       : in    std_logic;
          sample_f1_12       : in    std_logic;
          sample_f1_45       : in    std_logic;
          sample_f1_13       : in    std_logic;
          sample_f1_46       : in    std_logic;
          sample_f1_14       : in    std_logic;
          sample_f1_47       : in    std_logic;
          sample_f1_15       : in    std_logic;
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic;
          data_f1_out_valid  : out   std_logic;
          N_4                : in    std_logic;
          I_38_4             : in    std_logic;
          I_24_4             : in    std_logic;
          I_20_12            : in    std_logic;
          I_13_20            : in    std_logic;
          I_45_4             : in    std_logic;
          I_9_20             : in    std_logic;
          I_5_20             : in    std_logic;
          I_52_4             : in    std_logic;
          data_shaping_R1    : in    std_logic;
          data_shaping_R1_0  : in    std_logic;
          I_56_4             : in    std_logic;
          I_31_5             : in    std_logic;
          enable_f1          : in    std_logic;
          burst_f1           : in    std_logic;
          sample_f1_val_0    : in    std_logic;
          start_snapshot_f1  : in    std_logic
        );

end lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1;

architecture DEF_ARCH of 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_47_1, \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, 
        N_59, N_47_0, counter_points_snapshot_0_sqmuxa_1_0, 
        ADD_32x32_fast_I308_Y_0_0, 
        \counter_points_snapshot[28]_net_1\, 
        ADD_32x32_fast_I311_Y_0_0, 
        \counter_points_snapshot[31]_net_1\, 
        ADD_32x32_fast_I296_Y_0_0, 
        \un1_counter_points_snapshot[15]\, 
        ADD_32x32_fast_I310_Y_0_0, 
        \counter_points_snapshot[30]_net_1\, 
        ADD_32x32_fast_I309_Y_0_0, 
        \counter_points_snapshot[29]_net_1\, 
        ADD_32x32_fast_I304_Y_0_0, 
        \un1_counter_points_snapshot[7]\, 
        ADD_32x32_fast_I253_Y_0_0, N481, N485, 
        ADD_32x32_fast_I250_Y_2, ADD_32x32_fast_I250_Y_1, N483, 
        N487, N467, N470, N479, ADD_32x32_fast_I295_Y_0_0, 
        \counter_points_snapshot[15]_net_1\, 
        ADD_32x32_fast_I251_Y_2, ADD_32x32_fast_I251_Y_1, N489, 
        N464, ADD_32x32_fast_I302_Y_0_0, 
        \counter_points_snapshot[22]_net_1\, 
        ADD_32x32_fast_I252_Y_1, N550, ADD_32x32_fast_I294_Y_0_0, 
        \counter_points_snapshot[14]_net_1\, 
        ADD_32x32_fast_I303_Y_0_0, 
        \un1_counter_points_snapshot[8]\, 
        ADD_32x32_fast_I307_Y_0_0, 
        \un1_counter_points_snapshot[4]\, 
        ADD_32x32_fast_I301_Y_0_0, 
        \counter_points_snapshot[21]_net_1\, 
        ADD_32x32_fast_I288_Y_0_0, 
        \un1_counter_points_snapshot[23]\, 
        ADD_32x32_fast_I293_Y_0_0, 
        \counter_points_snapshot[13]_net_1\, 
        ADD_32x32_fast_I292_Y_0_0, 
        \un1_counter_points_snapshot[19]\, 
        ADD_32x32_fast_I300_Y_0_0, 
        \counter_points_snapshot[20]_net_1\, 
        ADD_32x32_fast_I306_Y_0_0, 
        \un1_counter_points_snapshot[5]\, 
        ADD_32x32_fast_I305_Y_0_0, 
        \un1_counter_points_snapshot[6]\, 
        ADD_32x32_fast_I299_Y_0_0, 
        \un1_counter_points_snapshot[12]\, 
        ADD_32x32_fast_I297_Y_0_0, 
        \un1_counter_points_snapshot[14]\, 
        ADD_32x32_fast_I254_Y_0, N554, ADD_32x32_fast_I298_Y_0_0, 
        \un1_counter_points_snapshot[13]\, 
        ADD_32x32_fast_I255_Y_0, N556, ADD_32x32_fast_I256_Y_0, 
        I112_un1_Y, N495, ADD_32x32_fast_I263_Y_0, N580, N588, 
        N533, ADD_32x32_fast_I282_Y_0_0, 
        \un1_counter_points_snapshot[29]\, 
        ADD_32x32_fast_I134_Y_1, N401, ADD_32x32_fast_I134_Y_0, 
        \un1_counter_points_snapshot[22]\, 
        \un1_counter_points_snapshot[25]\, 
        ADD_32x32_fast_I142_Y_0, 
        \un1_counter_points_snapshot[26]\, 
        \un1_counter_points_snapshot[27]\, 
        ADD_32x32_fast_I126_Y_1, 
        \un1_counter_points_snapshot[20]\, N419, 
        ADD_32x32_fast_I126_Y_0, 
        \un1_counter_points_snapshot[21]\, 
        ADD_32x32_fast_I118_Y_1, N425, ADD_32x32_fast_I118_Y_0, 
        N422, data_out_valid_9_i_0, un1_data_in_validlt30_27, 
        un1_data_in_validlt30_18, un1_data_in_validlt30_17, 
        un1_data_in_validlt30_23, un1_data_in_validlt30_26, 
        un1_data_in_validlt30_12, un1_data_in_validlt30_11, 
        un1_data_in_validlt30_22, un1_data_in_validlt30_25, 
        un1_data_in_validlt30_8, un1_data_in_validlt30_7, 
        un1_data_in_validlt30_20, un1_data_in_validlt30_2, 
        un1_data_in_validlt30_1, un1_data_in_validlt30_15, 
        un1_data_in_validlt30_14, 
        \counter_points_snapshot[27]_net_1\, 
        \counter_points_snapshot[26]_net_1\, 
        un1_data_in_validlt30_10, 
        \counter_points_snapshot[19]_net_1\, 
        \counter_points_snapshot[18]_net_1\, 
        un1_data_in_validlt30_6, 
        \counter_points_snapshot[11]_net_1\, 
        \counter_points_snapshot[10]_net_1\, 
        un1_data_in_validlt30_4, 
        \counter_points_snapshot[7]_net_1\, 
        \counter_points_snapshot[6]_net_1\, 
        \counter_points_snapshot[1]_net_1\, 
        \counter_points_snapshot[0]_net_1\, 
        \counter_points_snapshot[24]_net_1\, 
        \counter_points_snapshot[25]_net_1\, 
        \counter_points_snapshot[23]_net_1\, 
        \counter_points_snapshot[16]_net_1\, 
        \counter_points_snapshot[17]_net_1\, 
        \counter_points_snapshot[12]_net_1\, 
        \counter_points_snapshot[8]_net_1\, 
        \counter_points_snapshot[9]_net_1\, 
        \counter_points_snapshot[4]_net_1\, 
        \counter_points_snapshot[5]_net_1\, 
        \counter_points_snapshot[2]_net_1\, 
        \counter_points_snapshot[3]_net_1\, N758, N638, N622_i, 
        N654, N748, N628, N786, 
        \un1_data_out_valid_0_sqmuxa_2[10]\, 
        \un1_data_out_valid_0_sqmuxa_2[6]\, N652, 
        \un1_data_out_valid_0_sqmuxa_2[9]\, N789, N750_i, N630, 
        N744, N752, N_49, N_52, N_60, un1_data_in_validlto30_i, 
        N_47, counter_points_snapshot_0_sqmuxa_1, N740, N774, 
        N620, N738, N771_i, N618, 
        \un1_data_out_valid_0_sqmuxa_2[1]\, 
        \un1_counter_points_snapshot[30]\, N380, N756, N636, N529, 
        \un1_data_out_valid_0_sqmuxa_2[2]\, 
        \un1_data_out_valid_0_sqmuxa_2[8]\, N650, 
        \un1_data_out_valid_0_sqmuxa_2[4]\, N592, 
        \un1_data_out_valid_0_sqmuxa_2[3]\, 
        \un1_counter_points_snapshot[28]\, N594, 
        \un1_data_out_valid_0_sqmuxa_2[5]\, N766, N646, N443, 
        N440, N497, \un1_data_out_valid_0_sqmuxa_2[7]\, 
        \un1_counter_points_snapshot[24]\, N754, N634, N572, 
        \un1_data_out_valid_0_sqmuxa_2[11]\, N783, N742, N777, 
        N762, N642, N626, N764, N746, N574, N515, N511, N566, 
        N582, N_90, counter_points_snapshot_2_sqmuxa, N_94, 
        \counter_points_snapshot_10[6]\, 
        \counter_points_snapshot_10[10]\, N_25, N_35, 
        \sample_f1_wdata[32]\, \sample_f1_wdata[33]\, 
        \sample_f1_wdata[34]\, \sample_f1_wdata[35]\, 
        \sample_f1_wdata[19]\, \sample_f1_wdata[20]\, 
        \sample_f1_wdata[21]\, \sample_f1_wdata[22]\, 
        \sample_f1_wdata[23]\, \sample_f1_wdata[24]\, 
        \sample_f1_wdata[25]\, \sample_f1_wdata[26]\, 
        \sample_f1_wdata[27]\, \sample_f1_wdata[28]\, 
        \sample_f1_wdata[29]\, \sample_f1_wdata[30]\, 
        \sample_f1_wdata[31]\, \sample_f1_wdata[43]\, 
        \sample_f1_wdata[44]\, \sample_f1_wdata[45]\, 
        \sample_f1_wdata[46]\, \sample_f1_wdata[47]\, 
        \sample_f1_wdata[16]\, \sample_f1_wdata[17]\, 
        \sample_f1_wdata[18]\, \sample_f1_wdata[36]\, 
        \sample_f1_wdata[37]\, \sample_f1_wdata[38]\, 
        \sample_f1_wdata[39]\, \sample_f1_wdata[40]\, 
        \sample_f1_wdata[41]\, \sample_f1_wdata[42]\, N_9, N_7, 
        N780, N503, N570, N_27, \counter_points_snapshot_10[9]\, 
        N_93, N446, N_39, \counter_points_snapshot_10[1]\, N_85, 
        N_45, N_43, N_13, N_11, \counter_points_snapshot_10[2]\, 
        N_86, N_92, \counter_points_snapshot_10[8]\, N590, N531, 
        N527, N386, N383, \un1_counter_points_snapshot[31]\, 
        \un1_data_out_valid_0_sqmuxa_2[0]\, N_84, 
        \counter_points_snapshot_10[0]\, N586, N523, N_87, N_88, 
        \counter_points_snapshot_10[3]\, 
        \counter_points_snapshot_10[4]\, N_17, 
        \counter_points_snapshot_10[5]\, N_89, N519, N_31, N_29, 
        \counter_points_snapshot_10[7]\, N_91, N_33, N_41, 
        \counter_points_snapshot_10[11]\, N_95, N_21, N768, N_15, 
        N_37, N_23, N760, N_19, N578, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \counter_points_snapshot[13]\ : DFN1C0
      port map(D => N_9, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[13]_net_1\);
    
    \counter_points_snapshot[11]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[11]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[11]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I284_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[27]\, C => N592, Y => 
        \un1_data_out_valid_0_sqmuxa_2[4]\);
    
    \counter_points_snapshot_RNI7ND9[16]\ : NOR2
      port map(A => \counter_points_snapshot[16]_net_1\, B => 
        \counter_points_snapshot[17]_net_1\, Y => 
        un1_data_in_validlt30_8);
    
    \data_out[110]\ : DFN1C0
      port map(D => \sample_f1_wdata[46]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(110));
    
    \counter_points_snapshot_RNI9G66[8]\ : NOR2
      port map(A => \counter_points_snapshot[8]_net_1\, B => 
        \counter_points_snapshot[9]_net_1\, Y => 
        un1_data_in_validlt30_4);
    
    \counter_points_snapshot_RNO_0[10]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[10]\, B => 
        I_56_4, S => counter_points_snapshot_2_sqmuxa, Y => N_94);
    
    \counter_points_snapshot_RNO[27]\ : XA1C
      port map(A => N746, B => ADD_32x32_fast_I307_Y_0_0, C => 
        N_52, Y => N_37);
    
    \counter_points_snapshot[9]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[9]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[9]_net_1\);
    
    \counter_points_snapshot[28]\ : DFN1C0
      port map(D => N_39, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[28]_net_1\);
    
    \counter_points_snapshot_RNO[19]\ : XA1B
      port map(A => N762, B => ADD_32x32_fast_I299_Y_0_0, C => 
        N_52, Y => N_21);
    
    \data_out_RNO[96]\ : MX2
      port map(A => sample_f1_15, B => sample_f1_47, S => 
        data_shaping_R1_0, Y => \sample_f1_wdata[32]\);
    
    \data_out[91]\ : DFN1C0
      port map(D => \sample_f1_wdata[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(91));
    
    \counter_points_snapshot_RNISSL51[23]\ : NOR3C
      port map(A => un1_data_in_validlt30_12, B => 
        un1_data_in_validlt30_11, C => un1_data_in_validlt30_22, 
        Y => un1_data_in_validlt30_26);
    
    \data_out[120]\ : DFN1C0
      port map(D => sample_f1_wdata_56, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(120));
    
    \counter_points_snapshot_RNO[24]\ : XA1C
      port map(A => N752, B => ADD_32x32_fast_I304_Y_0_0, C => 
        N_52, Y => N_31);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y : OR3A
      port map(A => ADD_32x32_fast_I254_Y_0, B => N626, C => N783, 
        Y => N746);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I190_Y : NOR2
      port map(A => N586, B => N578, Y => N642);
    
    \data_out[130]\ : DFN1C0
      port map(D => sample_f1_wdata_66, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(130));
    
    \data_out[104]\ : DFN1C0
      port map(D => \sample_f1_wdata[40]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(104));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I104_Y : OR3B
      port map(A => N443, B => N446, C => N487, Y => N550);
    
    \counter_points_snapshot_RNO_0[4]\ : MX2C
      port map(A => I_20_12, B => 
        \un1_data_out_valid_0_sqmuxa_2[4]\, S => N_60, Y => N_88);
    
    \counter_points_snapshot_RNO_0[1]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[1]\, B => 
        I_5_20, S => counter_points_snapshot_2_sqmuxa, Y => N_85);
    
    \data_out[102]\ : DFN1C0
      port map(D => \sample_f1_wdata[38]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(102));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y : OR3B
      port map(A => N622_i, B => ADD_32x32_fast_I252_Y_1, C => 
        N777, Y => N742);
    
    \counter_points_snapshot_RNIHVMR1[11]\ : MX2
      port map(A => N_4, B => \counter_points_snapshot[11]_net_1\, 
        S => counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[20]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I282_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[29]\, B => 
        N_47_0, Y => ADD_32x32_fast_I282_Y_0_0);
    
    \counter_points_snapshot_RNO[7]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_91, Y => 
        \counter_points_snapshot_10[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I309_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I309_Y_0_0);
    
    \counter_points_snapshot_RNO[12]\ : XA1C
      port map(A => N780, B => ADD_32x32_fast_I292_Y_0_0, C => 
        N_52, Y => N_7);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I235_Y : NOR2
      port map(A => N650, B => N634, Y => N771_i);
    
    \data_out[93]\ : DFN1C0
      port map(D => \sample_f1_wdata[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(93));
    
    \counter_points_snapshot_RNIHME71[4]\ : MX2C
      port map(A => I_20_12, B => 
        \counter_points_snapshot[4]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[27]\);
    
    \counter_points_snapshot[4]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[4]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[4]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I301_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[21]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I301_Y_0_0);
    
    \data_out[159]\ : DFN1C0
      port map(D => sample_f1_wdata_95, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(159));
    
    \data_out[105]\ : DFN1C0
      port map(D => \sample_f1_wdata[41]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(105));
    
    \counter_points_snapshot[15]\ : DFN1C0
      port map(D => N_13, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[15]_net_1\);
    
    \data_out[141]\ : DFN1C0
      port map(D => sample_f1_wdata_77, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(141));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I108_Y : OR3B
      port map(A => N443, B => N446, C => N495, Y => N554);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I140_Y : OR2B
      port map(A => N527, B => N523, Y => N586);
    
    \data_out[81]\ : DFN1C0
      port map(D => \sample_f1_wdata[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(81));
    
    \counter_points_snapshot_RNIU5411[2]\ : MX2C
      port map(A => I_9_20, B => 
        \counter_points_snapshot[2]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[29]\);
    
    counter_points_snapshot_10_12_i_o2 : OR3B
      port map(A => enable_f1, B => N_60, C => burst_f1, Y => 
        N_52);
    
    \data_out_RNO[99]\ : MX2
      port map(A => sample_f1_12, B => sample_f1_44, S => 
        data_shaping_R1_0, Y => \sample_f1_wdata[35]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I310_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I310_Y_0_0);
    
    \data_out_RNO[104]\ : MX2
      port map(A => sample_f1_7, B => sample_f1_39, S => 
        data_shaping_R1, Y => \sample_f1_wdata[40]\);
    
    \counter_points_snapshot[7]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[7]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[7]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y_0 : OR3
      port map(A => I112_un1_Y, B => N495, C => N550, Y => 
        ADD_32x32_fast_I256_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I234_Y_0_o2 : 
        OR2A
      port map(A => N771_i, B => N425, Y => N768);
    
    \data_out[114]\ : DFN1C0
      port map(D => sample_f1_wdata_50, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(114));
    
    \counter_points_snapshot[0]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[0]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[0]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I182_Y : OR2
      port map(A => N578, B => N570, Y => N634);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I120_Y : NOR3
      port map(A => N419, B => N422, C => N503, Y => N566);
    
    \counter_points_snapshot[27]\ : DFN1C0
      port map(D => N_37, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[27]_net_1\);
    
    \data_out[143]\ : DFN1C0
      port map(D => sample_f1_wdata_79, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(143));
    
    \counter_points_snapshot_RNI319P[27]\ : NOR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[27]_net_1\, Y => 
        \un1_counter_points_snapshot[4]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I199_Y : OR2
      port map(A => N590, B => N533, Y => N654);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I110_Y : OR3C
      port map(A => N443, B => N440, C => N497, Y => N556);
    
    \data_out[112]\ : DFN1C0
      port map(D => sample_f1_wdata_48, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(112));
    
    \data_out[124]\ : DFN1C0
      port map(D => sample_f1_wdata_60, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(124));
    
    \data_out[134]\ : DFN1C0
      port map(D => sample_f1_wdata_70, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(134));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I80_Y : AO1
      port map(A => \un1_counter_points_snapshot[26]\, B => 
        \un1_counter_points_snapshot[25]\, C => N_47, Y => N523);
    
    \counter_points_snapshot_RNO[28]\ : XA1B
      port map(A => N744, B => ADD_32x32_fast_I308_Y_0_0, C => 
        N_52, Y => N_39);
    
    \data_out[83]\ : DFN1C0
      port map(D => \sample_f1_wdata[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(83));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_2 : NOR3A
      port map(A => ADD_32x32_fast_I250_Y_1, B => N483, C => N487, 
        Y => ADD_32x32_fast_I250_Y_2);
    
    \counter_points_snapshot_RNIMURI[26]\ : NOR3A
      port map(A => un1_data_in_validlt30_14, B => 
        \counter_points_snapshot[27]_net_1\, C => 
        \counter_points_snapshot[26]_net_1\, Y => 
        un1_data_in_validlt30_22);
    
    \data_out[122]\ : DFN1C0
      port map(D => sample_f1_wdata_58, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(122));
    
    \data_out[115]\ : DFN1C0
      port map(D => sample_f1_wdata_51, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(115));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I44_Y : OA1B
      port map(A => \un1_counter_points_snapshot[7]\, B => 
        \un1_counter_points_snapshot[8]\, C => N_47, Y => N487);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I38_Y_0_o2 : 
        OA1C
      port map(A => \un1_counter_points_snapshot[5]\, B => 
        \un1_counter_points_snapshot[4]\, C => N_47, Y => N481);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y_0 : AO1D
      port map(A => \un1_counter_points_snapshot[14]\, B => 
        N_47_1, C => N422, Y => ADD_32x32_fast_I118_Y_0);
    
    \data_out[132]\ : DFN1C0
      port map(D => sample_f1_wdata_68, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(132));
    
    \counter_points_snapshot_RNIM3VT[1]\ : MX2C
      port map(A => I_5_20, B => 
        \counter_points_snapshot[1]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[30]\);
    
    \counter_points_snapshot[30]\ : DFN1C0
      port map(D => N_43, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[30]_net_1\);
    
    \data_out[96]\ : DFN1C0
      port map(D => \sample_f1_wdata[32]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(96));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y : NOR3
      port map(A => N628, B => ADD_32x32_fast_I255_Y_0, C => N786, 
        Y => N748);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I294_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[14]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I294_Y_0_0);
    
    \data_out[125]\ : DFN1C0
      port map(D => sample_f1_wdata_61, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(125));
    
    \data_out[135]\ : DFN1C0
      port map(D => sample_f1_wdata_71, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(135));
    
    \data_out_RNO[87]\ : NOR2B
      port map(A => sample_f1_56, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[23]\);
    
    \data_out_RNO[108]\ : MX2
      port map(A => sample_f1_3, B => sample_f1_35, S => 
        data_shaping_R1, Y => \sample_f1_wdata[44]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I15_G0N : NOR3B
      port map(A => \counter_points_snapshot[15]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N425);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0 : NOR2
      port map(A => ADD_32x32_fast_I253_Y_0_0, B => N752, Y => 
        N744);
    
    data_out_valid : DFN1C0
      port map(D => N_49, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        data_f1_out_valid);
    
    \data_out_RNO[90]\ : NOR2B
      port map(A => sample_f1_53, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[26]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I174_Y : OR3
      port map(A => I112_un1_Y, B => N503, C => N570, Y => N626);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I29_G0N : OR3B
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N467);
    
    \data_out[71]\ : DFN1C0
      port map(D => sample_f1_wdata_7, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(71));
    
    \data_out[65]\ : DFN1C0
      port map(D => sample_f1_wdata_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(65));
    
    \counter_points_snapshot[18]\ : DFN1C0
      port map(D => N_19, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[18]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I260_Y : OR3B
      port map(A => N638, B => N622_i, C => N654, Y => N758);
    
    \data_out_RNO[98]\ : MX2
      port map(A => sample_f1_13, B => sample_f1_45, S => 
        data_shaping_R1_0, Y => \sample_f1_wdata[34]\);
    
    \data_out[86]\ : DFN1C0
      port map(D => \sample_f1_wdata[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(86));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I288_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[23]\, B => 
        N_47_0, Y => ADD_32x32_fast_I288_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I166_Y : OR3
      port map(A => I112_un1_Y, B => N503, C => N554, Y => N618);
    
    \data_out[150]\ : DFN1C0
      port map(D => sample_f1_wdata_86, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(150));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I297_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[14]\, B => 
        N_47_0, Y => ADD_32x32_fast_I297_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I296_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        N_47_0, Y => ADD_32x32_fast_I296_Y_0_0);
    
    \data_out[148]\ : DFN1C0
      port map(D => sample_f1_wdata_84, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(148));
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I13_G0N : NOR3B
      port map(A => \counter_points_snapshot[13]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N419);
    
    \counter_points_snapshot[8]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[8]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[8]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I178_Y : OR2A
      port map(A => N566, B => N574, Y => N630);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I136_Y : OR2B
      port map(A => N523, B => N519, Y => N582);
    
    \data_out[73]\ : DFN1C0
      port map(D => sample_f1_wdata_9, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(73));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \data_out[92]\ : DFN1C0
      port map(D => \sample_f1_wdata[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(92));
    
    \data_out[67]\ : DFN1C0
      port map(D => sample_f1_wdata_3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(67));
    
    \data_out[107]\ : DFN1C0
      port map(D => \sample_f1_wdata[43]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(107));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I14_G0N : NOR3B
      port map(A => \counter_points_snapshot[14]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N422);
    
    \counter_points_snapshot_RNISOQ14[6]\ : NOR3C
      port map(A => un1_data_in_validlt30_26, B => 
        un1_data_in_validlt30_25, C => un1_data_in_validlt30_27, 
        Y => un1_data_in_validlto30_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y_0 : OR3B
      port map(A => N580, B => N588, C => N533, Y => 
        ADD_32x32_fast_I263_Y_0);
    
    \counter_points_snapshot_RNO[6]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_90, Y => 
        \counter_points_snapshot_10[6]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I290_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[21]\, C => N786, Y => 
        \un1_data_out_valid_0_sqmuxa_2[10]\);
    
    \counter_points_snapshot[29]\ : DFN1C0
      port map(D => N_41, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[29]_net_1\);
    
    \data_out_RNO[94]\ : NOR2B
      port map(A => sample_f1_49, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[30]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I300_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I300_Y_0_0);
    
    \counter_points_snapshot_RNO[25]\ : XA1C
      port map(A => N750_i, B => ADD_32x32_fast_I305_Y_0_0, C => 
        N_52, Y => N_33);
    
    \counter_points_snapshot[20]\ : DFN1C0
      port map(D => N_23, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[20]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I302_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I302_Y_0_0);
    
    \counter_points_snapshot_RNI2T8P[26]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[26]_net_1\, Y => 
        \un1_counter_points_snapshot[5]\);
    
    \data_out_RNO[95]\ : NOR2B
      port map(A => sample_f1_48, B => data_shaping_R1, Y => 
        \sample_f1_wdata[31]\);
    
    \counter_points_snapshot[17]\ : DFN1C0
      port map(D => N_17, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[17]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I194_Y : OR2
      port map(A => N590, B => N582, Y => N646);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I88_Y : NOR2
      port map(A => N386, B => N383, Y => N531);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I292_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        N_47_0, Y => ADD_32x32_fast_I292_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I28_G0N : OR3B
      port map(A => \counter_points_snapshot[28]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N464);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y : OR3B
      port map(A => ADD_32x32_fast_I250_Y_2, B => N771_i, C => 
        N618, Y => N738);
    
    \data_out_RNO[93]\ : NOR2B
      port map(A => sample_f1_50, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[29]\);
    
    \data_out[154]\ : DFN1C0
      port map(D => sample_f1_wdata_90, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(154));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I261_Y_0_o2 : 
        OR2B
      port map(A => N764, B => N497, Y => N760);
    
    \data_out[82]\ : DFN1C0
      port map(D => \sample_f1_wdata[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(82));
    
    \data_out[117]\ : DFN1C0
      port map(D => sample_f1_wdata_53, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(117));
    
    \counter_points_snapshot_RNO[20]\ : XA1C
      port map(A => N760, B => ADD_32x32_fast_I300_Y_0_0, C => 
        N_52, Y => N_23);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y_0 : NOR3
      port map(A => N483, B => N487, C => N554, Y => 
        ADD_32x32_fast_I254_Y_0);
    
    \counter_points_snapshot_RNIICL51[14]\ : NOR3C
      port map(A => un1_data_in_validlt30_8, B => 
        un1_data_in_validlt30_7, C => un1_data_in_validlt30_20, Y
         => un1_data_in_validlt30_25);
    
    \data_out[76]\ : DFN1C0
      port map(D => sample_f1_wdata_12, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(76));
    
    \counter_points_snapshot_RNI1G66[4]\ : NOR2
      port map(A => \counter_points_snapshot[4]_net_1\, B => 
        \counter_points_snapshot[5]_net_1\, Y => 
        un1_data_in_validlt30_2);
    
    \data_out[152]\ : DFN1C0
      port map(D => sample_f1_wdata_88, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(152));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y_1 : AO1A
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[15]\, C => N425, Y => 
        ADD_32x32_fast_I118_Y_1);
    
    \counter_points_snapshot_RNIE0DC[6]\ : NOR3A
      port map(A => un1_data_in_validlt30_4, B => 
        \counter_points_snapshot[7]_net_1\, C => 
        \counter_points_snapshot[6]_net_1\, Y => 
        un1_data_in_validlt30_17);
    
    \data_out[149]\ : DFN1C0
      port map(D => sample_f1_wdata_85, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(149));
    
    \data_out[127]\ : DFN1C0
      port map(D => sample_f1_wdata_63, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(127));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I237_Y : OR2A
      port map(A => N638, B => N654, Y => N777);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I236_Y : NOR2
      port map(A => N652, B => N636, Y => N774);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I198_Y : OR2A
      port map(A => N588, B => N533, Y => N652);
    
    \data_out[137]\ : DFN1C0
      port map(D => sample_f1_wdata_73, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(137));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I30_G0N : OR3B
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N470);
    
    \data_out_RNO[81]\ : NOR2B
      port map(A => sample_f1_62, B => data_shaping_R1, Y => 
        \sample_f1_wdata[17]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I144_Y : OR2B
      port map(A => N531, B => N527, Y => N590);
    
    \data_out[155]\ : DFN1C0
      port map(D => sample_f1_wdata_91, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(155));
    
    \counter_points_snapshot_RNI1T8P[16]\ : NOR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[16]_net_1\, Y => 
        \un1_counter_points_snapshot[15]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \counter_points_snapshot_RNO[5]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_89, Y => 
        \counter_points_snapshot_10[5]\);
    
    \counter_points_snapshot_RNO[17]\ : XA1C
      port map(A => N766, B => ADD_32x32_fast_I297_Y_0_0, C => 
        N_52, Y => N_17);
    
    data_out_valid_RNO_0 : NOR2B
      port map(A => enable_f1, B => sample_f1_val_0, Y => 
        data_out_valid_9_i_0);
    
    \data_out[90]\ : DFN1C0
      port map(D => \sample_f1_wdata[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(90));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y_0 : AO1
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        \un1_counter_points_snapshot[21]\, C => N_47_1, Y => 
        ADD_32x32_fast_I126_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I124_Y : OR3
      port map(A => N419, B => N422, C => N511, Y => N570);
    
    \counter_points_snapshot[2]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[2]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[2]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y : OR3B
      port map(A => ADD_32x32_fast_I251_Y_2, B => N774, C => N620, 
        Y => N740);
    
    \counter_points_snapshot_RNO[14]\ : XA1C
      port map(A => N774, B => ADD_32x32_fast_I294_Y_0_0, C => 
        N_52, Y => N_11);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I20_G0N : OR3B
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N440);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I132_Y : OR2A
      port map(A => N519, B => N515, Y => N578);
    
    \counter_points_snapshot_RNI385K1[8]\ : MX2
      port map(A => I_45_4, B => 
        \counter_points_snapshot[8]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[23]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I282_Y_0 : XOR2
      port map(A => ADD_32x32_fast_I282_Y_0_0, B => N533, Y => 
        \un1_data_out_valid_0_sqmuxa_2[2]\);
    
    \data_out_RNO[92]\ : NOR2B
      port map(A => sample_f1_51, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[28]\);
    
    counter_points_snapshot_2_sqmuxa_0_a2 : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_60, Y => 
        counter_points_snapshot_2_sqmuxa);
    
    \data_out[99]\ : DFN1C0
      port map(D => \sample_f1_wdata[35]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(99));
    
    \counter_points_snapshot_RNI359P[18]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[18]_net_1\, Y => 
        \un1_counter_points_snapshot[13]\);
    
    \counter_points_snapshot_RNI219P[17]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[17]_net_1\, Y => 
        \un1_counter_points_snapshot[14]\);
    
    \data_out_RNO[100]\ : MX2
      port map(A => sample_f1_11, B => sample_f1_43, S => 
        data_shaping_R1, Y => \sample_f1_wdata[36]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I76_Y : OA1C
      port map(A => \un1_counter_points_snapshot[23]\, B => N_47, 
        C => N401, Y => N519);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I258_Y : NOR3
      port map(A => N634, B => N618, C => N650, Y => N754);
    
    \data_out[106]\ : DFN1C0
      port map(D => \sample_f1_wdata[42]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(106));
    
    \counter_points_snapshot_RNO[21]\ : XA1C
      port map(A => N758, B => ADD_32x32_fast_I301_Y_0_0, C => 
        N_52, Y => N_25);
    
    \data_out_RNO[103]\ : MX2
      port map(A => sample_f1_8, B => sample_f1_40, S => 
        data_shaping_R1, Y => \sample_f1_wdata[39]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I128_Y : OR2
      port map(A => N515, B => N511, Y => N574);
    
    \data_out[98]\ : DFN1C0
      port map(D => \sample_f1_wdata[34]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(98));
    
    \counter_points_snapshot_RNIEFFM1[6]\ : NOR3C
      port map(A => un1_data_in_validlt30_18, B => 
        un1_data_in_validlt30_17, C => un1_data_in_validlt30_23, 
        Y => un1_data_in_validlt30_27);
    
    \counter_points_snapshot_RNI1NC9[23]\ : NOR2
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        un1_data_in_validlt30_11);
    
    \data_out[80]\ : DFN1C0
      port map(D => \sample_f1_wdata[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(80));
    
    \data_out[72]\ : DFN1C0
      port map(D => sample_f1_wdata_8, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(72));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y : NOR3
      port map(A => N630, B => ADD_32x32_fast_I256_Y_0, C => N789, 
        Y => N750_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I22_G0N : OR3B
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N446);
    
    \counter_points_snapshot_RNITF66[2]\ : NOR2
      port map(A => \counter_points_snapshot[2]_net_1\, B => 
        \counter_points_snapshot[3]_net_1\, Y => 
        un1_data_in_validlt30_1);
    
    \counter_points_snapshot_RNI7C941[3]\ : MX2C
      port map(A => I_13_20, B => 
        \counter_points_snapshot[3]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[28]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I56_Y : AOI1
      port map(A => \un1_counter_points_snapshot[14]\, B => 
        \un1_counter_points_snapshot[13]\, C => N_47, Y => 
        I112_un1_Y);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I288_Y_0 : AX1B
      port map(A => N401, B => N650, C => 
        ADD_32x32_fast_I288_Y_0_0, Y => 
        \un1_data_out_valid_0_sqmuxa_2[8]\);
    
    \data_out_RNO[107]\ : MX2
      port map(A => sample_f1_4, B => sample_f1_36, S => 
        data_shaping_R1, Y => \sample_f1_wdata[43]\);
    
    counter_points_snapshot_2_sqmuxa_0_a2_0 : OR2A
      port map(A => start_snapshot_f1, B => sample_f1_val_0, Y
         => N_60);
    
    \data_out[89]\ : DFN1C0
      port map(D => \sample_f1_wdata[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(89));
    
    \counter_points_snapshot_RNIGRMR1[10]\ : MX2C
      port map(A => I_56_4, B => 
        \counter_points_snapshot[10]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[21]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y : NOR2
      port map(A => ADD_32x32_fast_I263_Y_0, B => N628, Y => N764);
    
    counter_points_snapshot_0_sqmuxa_1_0_a2 : OR3B
      port map(A => start_snapshot_f1, B => sample_f1_val_0, C
         => burst_f1, Y => counter_points_snapshot_0_sqmuxa_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I289_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[22]\, C => N789, Y => 
        \un1_data_out_valid_0_sqmuxa_2[9]\);
    
    \data_out_RNO[101]\ : MX2
      port map(A => sample_f1_10, B => sample_f1_42, S => 
        data_shaping_R1, Y => \sample_f1_wdata[37]\);
    
    \data_out[116]\ : DFN1C0
      port map(D => sample_f1_wdata_52, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(116));
    
    \counter_points_snapshot[19]\ : DFN1C0
      port map(D => N_21, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[19]_net_1\);
    
    \counter_points_snapshot_RNO_0[2]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[2]\, B => 
        I_9_20, S => counter_points_snapshot_2_sqmuxa, Y => N_86);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I298_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[13]\, B => 
        N_47_0, Y => ADD_32x32_fast_I298_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I197_Y : OR2
      port map(A => N594, B => N586, Y => N650);
    
    \counter_points_snapshot_RNI0L8P[24]\ : NOR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[24]_net_1\, Y => 
        \un1_counter_points_snapshot[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I285_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[26]\, C => N654, Y => 
        \un1_data_out_valid_0_sqmuxa_2[5]\);
    
    \counter_points_snapshot[10]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[10]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[10]_net_1\);
    
    \counter_points_snapshot_RNO[18]\ : XA1C
      port map(A => N764, B => ADD_32x32_fast_I298_Y_0_0, C => 
        N_52, Y => N_19);
    
    \data_out[88]\ : DFN1C0
      port map(D => \sample_f1_wdata[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(88));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_S_0 : XNOR2
      port map(A => \un1_counter_points_snapshot[31]\, B => N_47, 
        Y => \un1_data_out_valid_0_sqmuxa_2[0]\);
    
    \data_out[126]\ : DFN1C0
      port map(D => sample_f1_wdata_62, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(126));
    
    \data_out[94]\ : DFN1C0
      port map(D => \sample_f1_wdata[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(94));
    
    \data_out[140]\ : DFN1C0
      port map(D => sample_f1_wdata_76, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(140));
    
    \data_out[136]\ : DFN1C0
      port map(D => sample_f1_wdata_72, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(136));
    
    \counter_points_snapshot_RNI8HSA[0]\ : NOR3
      port map(A => \counter_points_snapshot[1]_net_1\, B => 
        \counter_points_snapshot[0]_net_1\, C => 
        \counter_points_snapshot[30]_net_1\, Y => 
        un1_data_in_validlt30_15);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I293_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[13]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I293_Y_0_0);
    
    \un1_data_out_valid_0_sqmuxa_1_i_0[31]\ : AOI1B
      port map(A => start_snapshot_f1, B => burst_f1, C => 
        sample_f1_val_0, Y => 
        \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\);
    
    \counter_points_snapshot_RNI8EQI[18]\ : NOR3A
      port map(A => un1_data_in_validlt30_10, B => 
        \counter_points_snapshot[19]_net_1\, C => 
        \counter_points_snapshot[18]_net_1\, Y => 
        un1_data_in_validlt30_20);
    
    \counter_points_snapshot_RNII6BN1[9]\ : MX2C
      port map(A => I_52_4, B => 
        \counter_points_snapshot[9]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[22]\);
    
    \counter_points_snapshot[22]\ : DFN1C0
      port map(D => N_27, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[22]_net_1\);
    
    \counter_points_snapshot_RNI57D9[24]\ : NOR2
      port map(A => \counter_points_snapshot[24]_net_1\, B => 
        \counter_points_snapshot[25]_net_1\, Y => 
        un1_data_in_validlt30_12);
    
    \data_out_RNO[86]\ : NOR2B
      port map(A => sample_f1_57, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[22]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I147_Y : OR2B
      port map(A => N531, B => N380, Y => N594);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I304_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[7]\, B => N_47_0, 
        Y => ADD_32x32_fast_I304_Y_0_0);
    
    \data_out[101]\ : DFN1C0
      port map(D => \sample_f1_wdata[37]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(101));
    
    \counter_points_snapshot_RNINKBE4[31]\ : OA1B
      port map(A => \counter_points_snapshot[31]_net_1\, B => 
        un1_data_in_validlto30_i, C => start_snapshot_f1, Y => 
        N_59);
    
    \data_out[157]\ : DFN1C0
      port map(D => sample_f1_wdata_93, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(157));
    
    \counter_points_snapshot_RNO[4]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_88, Y => 
        \counter_points_snapshot_10[4]\);
    
    \counter_points_snapshot_RNI37D9[14]\ : NOR2
      port map(A => \counter_points_snapshot[14]_net_1\, B => 
        \counter_points_snapshot[15]_net_1\, Y => 
        un1_data_in_validlt30_7);
    
    \counter_points_snapshot_RNO[30]\ : XA1C
      port map(A => N740, B => ADD_32x32_fast_I310_Y_0_0, C => 
        N_52, Y => N_43);
    
    \counter_points_snapshot[6]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[6]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[6]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I54_Y_0_o2 : AO1
      port map(A => \un1_counter_points_snapshot[13]\, B => 
        \un1_counter_points_snapshot[12]\, C => N_47, Y => N497);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I176_Y : OR3
      port map(A => ADD_32x32_fast_I118_Y_0, B => 
        ADD_32x32_fast_I118_Y_1, C => N572, Y => N628);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y_0 : AOI1
      port map(A => \un1_counter_points_snapshot[22]\, B => 
        \un1_counter_points_snapshot[25]\, C => N_47_1, Y => 
        ADD_32x32_fast_I134_Y_0);
    
    \data_out[70]\ : DFN1C0
      port map(D => sample_f1_wdata_6, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(70));
    
    \counter_points_snapshot_RNO_0[5]\ : MX2C
      port map(A => I_24_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[5]\, S => N_60, Y => N_89);
    
    \data_out[84]\ : DFN1C0
      port map(D => \sample_f1_wdata[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(84));
    
    \data_out[103]\ : DFN1C0
      port map(D => \sample_f1_wdata[39]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(103));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I7_G0N : NOR2
      port map(A => \un1_counter_points_snapshot[24]\, B => N_47, 
        Y => N401);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I84_Y : AO1
      port map(A => \un1_counter_points_snapshot[28]\, B => 
        \un1_counter_points_snapshot[27]\, C => N_47, Y => N527);
    
    \counter_points_snapshot[5]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[5]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[5]_net_1\);
    
    \counter_points_snapshot_RNO[26]\ : XA1C
      port map(A => N748, B => ADD_32x32_fast_I306_Y_0_0, C => 
        N_52, Y => N_35);
    
    \data_out[79]\ : DFN1C0
      port map(D => sample_f1_wdata_15, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(79));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I281_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[30]\, C => N380, Y => 
        \un1_data_out_valid_0_sqmuxa_2[1]\);
    
    \counter_points_snapshot_RNITC8P[12]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1_0, B => 
        \counter_points_snapshot[12]_net_1\, Y => 
        \un1_counter_points_snapshot[19]\);
    
    \data_out[144]\ : DFN1C0
      port map(D => sample_f1_wdata_80, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(144));
    
    counter_points_snapshot_0_sqmuxa_1_0_a2_0 : OR3B
      port map(A => start_snapshot_f1, B => sample_f1_val_0, C
         => burst_f1, Y => counter_points_snapshot_0_sqmuxa_1_0);
    
    \data_out_RNO[89]\ : NOR2B
      port map(A => sample_f1_54, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[25]\);
    
    \counter_points_snapshot_RNO[8]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_92, Y => 
        \counter_points_snapshot_10[8]\);
    
    \data_out[111]\ : DFN1C0
      port map(D => \sample_f1_wdata[47]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(111));
    
    \counter_points_snapshot_RNID7E9[28]\ : NOR2
      port map(A => \counter_points_snapshot[28]_net_1\, B => 
        \counter_points_snapshot[29]_net_1\, Y => 
        un1_data_in_validlt30_14);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I295_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[15]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I295_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_CO1 : OR2A
      port map(A => \un1_counter_points_snapshot[31]\, B => 
        N_47_1, Y => N380);
    
    \data_out[142]\ : DFN1C0
      port map(D => sample_f1_wdata_78, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(142));
    
    \data_out[78]\ : DFN1C0
      port map(D => sample_f1_wdata_14, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(78));
    
    \counter_points_snapshot_RNO[23]\ : XA1B
      port map(A => N754, B => ADD_32x32_fast_I303_Y_0_0, C => 
        N_52, Y => N_29);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I184_Y : OR2A
      port map(A => N580, B => N572, Y => N636);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y_1 : AO1A
      port map(A => N_47_0, B => 
        \un1_counter_points_snapshot[23]\, C => N401, Y => 
        ADD_32x32_fast_I134_Y_1);
    
    \counter_points_snapshot_RNO_0[3]\ : MX2C
      port map(A => I_13_20, B => 
        \un1_data_out_valid_0_sqmuxa_2[3]\, S => N_60, Y => N_87);
    
    \counter_points_snapshot[26]\ : DFN1C0
      port map(D => N_35, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[26]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I305_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[6]\, B => N_47_0, 
        Y => ADD_32x32_fast_I305_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y_1 : NOR3
      port map(A => N479, B => N483, C => N550, Y => 
        ADD_32x32_fast_I252_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I1_G0N : NOR2
      port map(A => \un1_counter_points_snapshot[30]\, B => 
        N_47_1, Y => N383);
    
    \data_out[121]\ : DFN1C0
      port map(D => sample_f1_wdata_57, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(121));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I60_Y : AO1A
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[15]\, C => N425, Y => N503);
    
    \counter_points_snapshot_RNO[0]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_84, Y => 
        \counter_points_snapshot_10[0]\);
    
    \data_out[131]\ : DFN1C0
      port map(D => sample_f1_wdata_67, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(131));
    
    \data_out[113]\ : DFN1C0
      port map(D => sample_f1_wdata_49, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(113));
    
    \counter_points_snapshot_RNIS4KA1[5]\ : MX2C
      port map(A => I_24_4, B => 
        \counter_points_snapshot[5]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[26]\);
    
    \data_out[145]\ : DFN1C0
      port map(D => sample_f1_wdata_81, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(145));
    
    \data_out[66]\ : DFN1C0
      port map(D => sample_f1_wdata_2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(66));
    
    \counter_points_snapshot[1]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[1]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[1]_net_1\);
    
    \counter_points_snapshot_RNO[31]\ : XA1B
      port map(A => N738, B => ADD_32x32_fast_I311_Y_0_0, C => 
        N_52, Y => N_45);
    
    \data_out_RNO[109]\ : MX2
      port map(A => sample_f1_2, B => sample_f1_34, S => 
        data_shaping_R1, Y => \sample_f1_wdata[45]\);
    
    \counter_points_snapshot_RNO_0[0]\ : MX2B
      port map(A => nb_snapshot_param(0), B => 
        \un1_data_out_valid_0_sqmuxa_2[0]\, S => N_60, Y => N_84);
    
    \counter_points_snapshot_RNO[15]\ : XA1C
      port map(A => N771_i, B => ADD_32x32_fast_I295_Y_0_0, C => 
        N_52, Y => N_13);
    
    \data_out[123]\ : DFN1C0
      port map(D => sample_f1_wdata_59, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(123));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \counter_points_snapshot_RNILDVG1[7]\ : MX2C
      port map(A => I_38_4, B => 
        \counter_points_snapshot[7]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[24]\);
    
    \data_out[133]\ : DFN1C0
      port map(D => sample_f1_wdata_69, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(133));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I21_G0N : OR3B
      port map(A => \counter_points_snapshot[21]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N443);
    
    \counter_points_snapshot_RNO[29]\ : XA1C
      port map(A => N742, B => ADD_32x32_fast_I309_Y_0_0, C => 
        N_52, Y => N_41);
    
    \counter_points_snapshot_RNI5OT25_1[31]\ : OR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, 
        B => N_59, Y => N_47);
    
    \counter_points_snapshot[31]\ : DFN1C0
      port map(D => N_45, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[31]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I36_Y : AO1C
      port map(A => N_47, B => \un1_counter_points_snapshot[4]\, 
        C => N464, Y => N479);
    
    \counter_points_snapshot_RNI1P8P[25]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[25]_net_1\, Y => 
        \un1_counter_points_snapshot[6]\);
    
    \data_out_RNO[97]\ : MX2
      port map(A => sample_f1_14, B => sample_f1_46, S => 
        data_shaping_R1_0, Y => \sample_f1_wdata[33]\);
    
    \data_out[74]\ : DFN1C0
      port map(D => sample_f1_wdata_10, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(74));
    
    \counter_points_snapshot_RNO[10]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_94, Y => 
        \counter_points_snapshot_10[10]\);
    
    \data_out[108]\ : DFN1C0
      port map(D => \sample_f1_wdata[44]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(108));
    
    \counter_points_snapshot_RNO_0[6]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[6]\, B => 
        I_31_5, S => counter_points_snapshot_2_sqmuxa, Y => N_90);
    
    \counter_points_snapshot_RNIF5QQ[0]\ : MX2A
      port map(A => nb_snapshot_param(0), B => 
        \counter_points_snapshot[0]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[31]\);
    
    \data_out[156]\ : DFN1C0
      port map(D => sample_f1_wdata_92, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(156));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I240_Y : OR3B
      port map(A => N580, B => N588, C => N533, Y => N786);
    
    \data_out_RNO[106]\ : MX2
      port map(A => sample_f1_5, B => sample_f1_37, S => 
        data_shaping_R1, Y => \sample_f1_wdata[42]\);
    
    \counter_points_snapshot_RNO_0[8]\ : MX2C
      port map(A => I_45_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[8]\, S => N_60, Y => N_92);
    
    \data_out_RNO[80]\ : NOR2B
      port map(A => sample_f1_63, B => data_shaping_R1, Y => 
        \sample_f1_wdata[16]\);
    
    \counter_points_snapshot_RNO[1]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_85, Y => 
        \counter_points_snapshot_10[1]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I303_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[8]\, B => N_47_0, 
        Y => ADD_32x32_fast_I303_Y_0_0);
    
    \counter_points_snapshot_RNIT6C9[20]\ : NOR2
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        \counter_points_snapshot[21]_net_1\, Y => 
        un1_data_in_validlt30_10);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I40_Y : AOI1
      port map(A => \un1_counter_points_snapshot[6]\, B => 
        \un1_counter_points_snapshot[5]\, C => N_47, Y => N483);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I257_Y_0_o2 : 
        OR2
      port map(A => N756, B => N489, Y => N752);
    
    \counter_points_snapshot_RNO[22]\ : XA1C
      port map(A => N756, B => ADD_32x32_fast_I302_Y_0_0, C => 
        N_52, Y => N_27);
    
    \data_out_RNO[88]\ : NOR2B
      port map(A => sample_f1_55, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[24]\);
    
    \counter_points_snapshot_RNIQTOI[10]\ : NOR3A
      port map(A => un1_data_in_validlt30_6, B => 
        \counter_points_snapshot[11]_net_1\, C => 
        \counter_points_snapshot[10]_net_1\, Y => 
        un1_data_in_validlt30_18);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I146_Y : NOR2
      port map(A => N533, B => N529, Y => N592);
    
    \counter_points_snapshot[12]\ : DFN1C0
      port map(D => N_7, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[12]_net_1\);
    
    \counter_points_snapshot[24]\ : DFN1C0
      port map(D => N_31, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[24]_net_1\);
    
    \counter_points_snapshot_RNI6H9N[0]\ : NOR3C
      port map(A => un1_data_in_validlt30_2, B => 
        un1_data_in_validlt30_1, C => un1_data_in_validlt30_15, Y
         => un1_data_in_validlt30_23);
    
    \data_out[95]\ : DFN1C0
      port map(D => \sample_f1_wdata[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(95));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y : OR2B
      port map(A => ADD_32x32_fast_I126_Y_1, B => 
        ADD_32x32_fast_I126_Y_0, Y => N572);
    
    \data_out_RNO[110]\ : MX2
      port map(A => sample_f1_1, B => sample_f1_33, S => 
        data_shaping_R1, Y => \sample_f1_wdata[46]\);
    
    \counter_points_snapshot_RNIVMC9[12]\ : NOR2
      port map(A => \counter_points_snapshot[12]_net_1\, B => 
        \counter_points_snapshot[13]_net_1\, Y => 
        un1_data_in_validlt30_6);
    
    \counter_points_snapshot_RNO_0[9]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[9]\, B => 
        I_52_4, S => counter_points_snapshot_2_sqmuxa, Y => N_93);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y_1 : OA1C
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        N_47_1, C => N419, Y => ADD_32x32_fast_I126_Y_1);
    
    \counter_points_snapshot_RNO[3]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_87, Y => 
        \counter_points_snapshot_10[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y_0 : AOI1
      port map(A => \un1_counter_points_snapshot[26]\, B => 
        \un1_counter_points_snapshot[27]\, C => N_47_1, Y => 
        ADD_32x32_fast_I142_Y_0);
    
    \data_out[118]\ : DFN1C0
      port map(D => sample_f1_wdata_54, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(118));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I241_Y : OR2A
      port map(A => N380, B => N646, Y => N789);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I306_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[5]\, B => N_47_0, 
        Y => ADD_32x32_fast_I306_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_1 : NOR3B
      port map(A => N467, B => N464, C => N481, Y => 
        ADD_32x32_fast_I251_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I239_Y : OR2A
      port map(A => N642, B => N594, Y => N783);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I287_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[24]\, C => N650, Y => 
        \un1_data_out_valid_0_sqmuxa_2[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I286_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[25]\, C => N652, Y => 
        \un1_data_out_valid_0_sqmuxa_2[6]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I46_Y_0_o2 : 
        AO1C
      port map(A => N_47, B => \un1_counter_points_snapshot[8]\, 
        C => N446, Y => N489);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I291_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[20]\, C => N783, Y => 
        \un1_data_out_valid_0_sqmuxa_2[11]\);
    
    \data_out[128]\ : DFN1C0
      port map(D => sample_f1_wdata_64, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(128));
    
    \counter_points_snapshot_RNO[11]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_95, Y => 
        \counter_points_snapshot_10[11]\);
    
    \data_out[97]\ : DFN1C0
      port map(D => \sample_f1_wdata[33]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(97));
    
    \data_out[138]\ : DFN1C0
      port map(D => sample_f1_wdata_74, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(138));
    
    \data_out_RNO[84]\ : NOR2B
      port map(A => sample_f1_59, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[20]\);
    
    \data_out[85]\ : DFN1C0
      port map(D => \sample_f1_wdata[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(85));
    
    \counter_points_snapshot[3]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[3]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[3]_net_1\);
    
    \data_out_RNO[85]\ : NOR2B
      port map(A => sample_f1_58, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[21]\);
    
    \data_out[109]\ : DFN1C0
      port map(D => \sample_f1_wdata[45]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(109));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I68_Y : OA1C
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        \un1_counter_points_snapshot[20]\, C => N_47, Y => N511);
    
    \data_out_RNO[111]\ : MX2
      port map(A => sample_f1_0, B => sample_f1_32, S => 
        data_shaping_R1, Y => \sample_f1_wdata[47]\);
    
    \counter_points_snapshot[23]\ : DFN1C0
      port map(D => N_29, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[23]_net_1\);
    
    \counter_points_snapshot[21]\ : DFN1C0
      port map(D => N_25, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[21]_net_1\);
    
    \counter_points_snapshot[16]\ : DFN1C0
      port map(D => N_15, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[16]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y_0 : OR3
      port map(A => N485, B => N489, C => N556, Y => 
        ADD_32x32_fast_I255_Y_0);
    
    \data_out[147]\ : DFN1C0
      port map(D => sample_f1_wdata_83, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(147));
    
    \data_out[151]\ : DFN1C0
      port map(D => sample_f1_wdata_87, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(151));
    
    \data_out_RNO[83]\ : NOR2B
      port map(A => sample_f1_60, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[19]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I299_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[12]\, B => 
        N_47_0, Y => ADD_32x32_fast_I299_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I308_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[28]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I308_Y_0_0);
    
    \data_out[87]\ : DFN1C0
      port map(D => \sample_f1_wdata[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(87));
    
    \data_out[153]\ : DFN1C0
      port map(D => sample_f1_wdata_89, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(153));
    
    \counter_points_snapshot_RNI499P[19]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[19]_net_1\, Y => 
        \un1_counter_points_snapshot[12]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I283_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[28]\, C => N594, Y => 
        \un1_data_out_valid_0_sqmuxa_2[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I259_Y : OR3
      port map(A => N636, B => N620, C => N652, Y => N756);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I86_Y : AO1D
      port map(A => \un1_counter_points_snapshot[28]\, B => N_47, 
        C => N386, Y => N529);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y : NOR2
      port map(A => ADD_32x32_fast_I142_Y_0, B => N529, Y => N588);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I307_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[4]\, B => N_47_0, 
        Y => ADD_32x32_fast_I307_Y_0_0);
    
    \data_out_RNO[91]\ : NOR2B
      port map(A => sample_f1_52, B => data_shaping_R1_0, Y => 
        \sample_f1_wdata[27]\);
    
    \data_out[119]\ : DFN1C0
      port map(D => sample_f1_wdata_55, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(119));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_1 : NOR3B
      port map(A => N467, B => N470, C => N479, Y => 
        ADD_32x32_fast_I250_Y_1);
    
    \counter_points_snapshot_RNI5OT25[31]\ : OR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, 
        B => N_59, Y => N_47_1);
    
    \data_out_RNO[102]\ : MX2
      port map(A => sample_f1_9, B => sample_f1_41, S => 
        data_shaping_R1, Y => \sample_f1_wdata[38]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I72_Y : AOI1
      port map(A => \un1_counter_points_snapshot[22]\, B => 
        \un1_counter_points_snapshot[21]\, C => N_47, Y => N515);
    
    \counter_points_snapshot_RNO_0[7]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[7]\, B => 
        I_38_4, S => counter_points_snapshot_2_sqmuxa, Y => N_91);
    
    \counter_points_snapshot_RNO[9]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_93, Y => 
        \counter_points_snapshot_10[9]\);
    
    \counter_points_snapshot_RNI5OT25_0[31]\ : OR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, 
        B => N_59, Y => N_47_0);
    
    \data_out[69]\ : DFN1C0
      port map(D => sample_f1_wdata_5, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(69));
    
    \data_out[129]\ : DFN1C0
      port map(D => sample_f1_wdata_65, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(129));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I311_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[31]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I311_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_2 : NOR3A
      port map(A => ADD_32x32_fast_I251_Y_1, B => N485, C => N489, 
        Y => ADD_32x32_fast_I251_Y_2);
    
    \data_out[139]\ : DFN1C0
      port map(D => sample_f1_wdata_75, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(139));
    
    \counter_points_snapshot[25]\ : DFN1C0
      port map(D => N_33, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[25]_net_1\);
    
    \data_out_RNO[82]\ : NOR2B
      port map(A => sample_f1_61, B => data_shaping_R1, Y => 
        \sample_f1_wdata[18]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y : NOR2
      port map(A => ADD_32x32_fast_I134_Y_1, B => 
        ADD_32x32_fast_I134_Y_0, Y => N580);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I238_Y_0_o2 : 
        OA1C
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        N_47_1, C => N783, Y => N780);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I90_Y : OR2A
      port map(A => N380, B => N383, Y => N533);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I42_Y : OA1C
      port map(A => \un1_counter_points_snapshot[6]\, B => 
        \un1_counter_points_snapshot[7]\, C => N_47, Y => N485);
    
    \data_out[75]\ : DFN1C0
      port map(D => sample_f1_wdata_11, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(75));
    
    \data_out[68]\ : DFN1C0
      port map(D => sample_f1_wdata_4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(68));
    
    \counter_points_snapshot_RNO_0[11]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[11]\, B => N_4, 
        S => counter_points_snapshot_2_sqmuxa, Y => N_95);
    
    \counter_points_snapshot[14]\ : DFN1C0
      port map(D => N_11, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[14]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I52_Y : OAI1
      port map(A => N_47, B => \un1_counter_points_snapshot[12]\, 
        C => N440, Y => N495);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I168_Y : OR3
      port map(A => ADD_32x32_fast_I118_Y_0, B => 
        ADD_32x32_fast_I118_Y_1, C => N556, Y => N620);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I264_Y : NOR3A
      port map(A => N380, B => N646, C => N630, Y => N766);
    
    \counter_points_snapshot_RNIVG8P[23]\ : NOR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        \un1_counter_points_snapshot[8]\);
    
    \counter_points_snapshot_RNO[16]\ : XA1C
      port map(A => N768, B => ADD_32x32_fast_I296_Y_0_0, C => 
        N_52, Y => N_15);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I170_Y : NOR3A
      port map(A => N566, B => I112_un1_Y, C => N495, Y => N622_i);
    
    \counter_points_snapshot_RNI8NPD1[6]\ : MX2C
      port map(A => I_31_5, B => 
        \counter_points_snapshot[6]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[25]\);
    
    data_out_valid_RNO : OA1A
      port map(A => N_59, B => burst_f1, C => 
        data_out_valid_9_i_0, Y => N_49);
    
    \data_out[100]\ : DFN1C0
      port map(D => \sample_f1_wdata[36]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(100));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I262_Y : OR3A
      port map(A => N642, B => N594, C => N626, Y => N762);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0_0 : OR2
      port map(A => N481, B => N485, Y => 
        ADD_32x32_fast_I253_Y_0_0);
    
    \data_out[77]\ : DFN1C0
      port map(D => sample_f1_wdata_13, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(77));
    
    \data_out[146]\ : DFN1C0
      port map(D => sample_f1_wdata_82, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(146));
    
    \counter_points_snapshot_RNO[2]\ : NOR3A
      port map(A => enable_f1, B => burst_f1, C => N_86, Y => 
        \counter_points_snapshot_10[2]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I186_Y : NOR2
      port map(A => N582, B => N574, Y => N638);
    
    \counter_points_snapshot_RNO[13]\ : XA1B
      port map(A => N777, B => ADD_32x32_fast_I293_Y_0_0, C => 
        N_52, Y => N_9);
    
    \data_out[158]\ : DFN1C0
      port map(D => sample_f1_wdata_94, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(158));
    
    \data_out_RNO[105]\ : MX2
      port map(A => sample_f1_6, B => sample_f1_38, S => 
        data_shaping_R1, Y => \sample_f1_wdata[41]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I2_G0N : NOR2
      port map(A => \un1_counter_points_snapshot[29]\, B => N_47, 
        Y => N386);
    
    \data_out[64]\ : DFN1C0
      port map(D => sample_f1_wdata_0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f1_out(64));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_snapshot_controler is

    port( delta_f2_f0       : in    std_logic_vector(9 downto 0);
          delta_snapshot    : in    std_logic_vector(15 downto 0);
          delta_f2_f1       : in    std_logic_vector(9 downto 0);
          start_snapshot_f2 : out   std_logic;
          start_snapshot_f1 : out   std_logic;
          start_snapshot_f0 : out   std_logic;
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          sample_f0_val_0   : in    std_logic;
          sample_f2_val     : in    std_logic;
          coarse_time_0_c   : in    std_logic
        );

end lpp_waveform_snapshot_controler;

architecture DEF_ARCH of lpp_waveform_snapshot_controler is 

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AXOI2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_34, N_80, \counter_delta_f0[26]_net_1\, N_57_0, 
        N_265, \counter_delta_f0[19]_net_1\, N_105, 
        counter_delta_f0_n19, N_106, N_57, counter_delta_f0_n20, 
        \counter_delta_f0[20]_net_1\, N_89, 
        \counter_delta_f0[0]_net_1\, \counter_delta_f0[1]_net_1\, 
        \counter_delta_f0[2]_net_1\, N_99, N_67, 
        \counter_delta_f0[11]_net_1\, 
        \counter_delta_f0[12]_net_1\, N_101, 
        \counter_delta_f0[13]_net_1\, 
        \counter_delta_f0[14]_net_1\, N_103, 
        \counter_delta_f0[15]_net_1\, 
        \counter_delta_f0[16]_net_1\, 
        \counter_delta_f0[17]_net_1\, 
        \counter_delta_f0[18]_net_1\, N_276, N_58, 
        \counter_delta_f0[21]_net_1\, N_277, N_86_i, N_28, N_62, 
        \counter_delta_f0[23]_net_1\, N_30, N_98_i, N_32, N_66, 
        \counter_delta_f0[25]_net_1\, 
        \counter_delta_f0[22]_net_1\, 
        \counter_delta_f0[24]_net_1\, N_63, 
        \counter_delta_f0[9]_net_1\, \counter_delta_f0[10]_net_1\, 
        N_59, \counter_delta_f0[7]_net_1\, 
        \counter_delta_f0[8]_net_1\, N_55, 
        \counter_delta_f0[5]_net_1\, \counter_delta_f0[6]_net_1\, 
        \counter_delta_f0[3]_net_1\, \counter_delta_f0[4]_net_1\, 
        un2_coarse_time_0_0, \coarse_time_0_r\, N_504_0, 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, N_9_0, 
        N_9_tz, N_7, \start_snapshot_fothers_temp\, 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, 
        \counter_delta_snapshot_e27_0_0_o2_m6_e_3\, 
        counter_delta_snapshot_e27_0_0_o2_m6_e_2, N_398, 
        start_snapshot_f22_0_a2_11_0_a2_3_i, 
        \counter_delta_snapshot[23]_net_1\, 
        \counter_delta_snapshot[22]_net_1\, 
        start_snapshot_f22_0_a2_11_0_a2_2_i, 
        \counter_delta_snapshot[19]_net_1\, 
        \counter_delta_snapshot[18]_net_1\, N_495, 
        \counter_delta_snapshot[12]_net_1\, 
        start_snapshot_f2_temp3_0_a2_0, start_snapshot_f22_11_i, 
        start_snapshot_f22_10, start_snapshot_f22_0_a2_1, 
        start_snapshot_f22_0_a2_0, 
        start_snapshot_f22_0_a2_11_0_a2_2_0, 
        un12_start_snapshot_fothers_temp_NE, 
        un12_start_snapshot_fothers_temp_NE_12, 
        un12_start_snapshot_fothers_temp_NE_13, N_493, 
        \counter_delta_snapshot_e12_i_0_a2_0\, 
        start_snapshot_f2_temp3, counter_delta_snapshot_e12_i_0_0, 
        counter_delta_snapshot_e25_0_0_0, 
        \counter_delta_snapshot[25]_net_1\, N_421, 
        counter_delta_snapshot_e25_0_0_a2_0, 
        counter_delta_snapshot_e23_0_0_0, N_189, 
        counter_delta_snapshot_e8_i_0, 
        counter_delta_snapshot_e8_i_a2_0, N_466, 
        counter_delta_snapshot_e2_i_0, 
        counter_delta_snapshot_e2_i_a2_0, N_436, 
        counter_delta_snapshot_e3_i_0, 
        \counter_delta_snapshot[3]_net_1\, N_440, 
        counter_delta_snapshot_e6_i_0, 
        \counter_delta_snapshot[6]_net_1\, N_455, 
        counter_delta_snapshot_e7_i_0, 
        \counter_delta_snapshot[7]_net_1\, N_460, 
        counter_delta_snapshot_e9_i_0, 
        counter_delta_snapshot_e9_i_a2_0, N_470, 
        counter_delta_snapshot_e15_i_0_0, 
        \counter_delta_snapshot[15]_net_1\, N_478, 
        counter_delta_snapshot_e14_i_0_0, 
        \counter_delta_snapshot[14]_net_1\, N_484, 
        counter_delta_snapshot_e13_i_0_0, 
        \counter_delta_snapshot[13]_net_1\, N_285, 
        counter_delta_snapshot_e4_i_0, 
        \counter_delta_snapshot[4]_net_1\, N_445, 
        counter_delta_snapshot_e5_i_0, 
        \counter_delta_snapshot_i[5]\, N_450, 
        counter_delta_snapshot_e11_i_0_0, 
        counter_delta_snapshot_e11_i_0_a2_0, N_294, 
        counter_delta_snapshot_e0_i_0, 
        \counter_delta_snapshot[0]_net_1\, 
        counter_delta_snapshot_e10_i_0, 
        \counter_delta_snapshot[10]_net_1\, N_474, 
        counter_delta_f0_n18_0_0_a2_0, 
        counter_delta_snapshot_e16_i_i_0, 
        \counter_delta_snapshot[16]_net_1\, N_168, 
        counter_delta_snapshot_e19_i_i_0, 
        counter_delta_snapshot_e19_i_i_a2_0, N_178, 
        counter_delta_snapshot_e21_0_0_0, 
        \counter_delta_snapshot[21]_net_1\, un2_coarse_time_0, 
        N_183, counter_delta_snapshot_e13_i_0_a2_2_0, N_393, 
        counter_delta_snapshot_e23_0_0_a2_0, 
        counter_delta_f0_n16_0_0_a2_0, 
        counter_delta_snapshot_e21_0_0_a2_0, 
        \counter_delta_snapshot_RNI0DDG1[7]_net_1\, 
        \counter_delta_snapshot[8]_net_1\, N_388, 
        \counter_delta_snapshot[2]_net_1\, N_382, 
        counter_delta_snapshot_e6_i_a2_0, N_386, 
        counter_delta_snapshot_e7_i_a2_0, N_387, 
        \counter_delta_snapshot[9]_net_1\, N_389, 
        counter_delta_snapshot_e15_i_0_a2_0, N_395, 
        counter_delta_snapshot_e14_i_0_a2_0, N_394, 
        counter_delta_snapshot_e13_i_0_a2_0, 
        counter_delta_snapshot_e16_i_i_a2_0, N_396, 
        counter_delta_snapshot_e4_i_a2_0, N_384, 
        counter_delta_snapshot_e5_i_a2_0, N_385, 
        \counter_delta_snapshot_i[11]\, N_391, 
        counter_delta_f0_n14_0_0_a2_0, 
        \counter_delta_snapshot_e27_0_0_o2_m6_e_1\, 
        start_snapshot_f22_0_a2_11_0_a2_1, 
        \counter_delta_snapshot[26]_net_1\, 
        \counter_delta_snapshot[24]_net_1\, 
        counter_delta_f0_n12_0_0_a2_0, counter_delta_f0_n10_0_i_0, 
        counter_delta_f0lde_i_a2_0_1_3, 
        counter_delta_f0lde_i_a2_0_1_2, counter_delta_f0_1_0_a2_7, 
        N_273, counter_delta_f0_1_0_a2_2_0, 
        start_snapshot_f12_0_a2_7, start_snapshot_f12_0_a2_1, 
        start_snapshot_f12_0_a2_0, start_snapshot_f12_0_a2_4, 
        start_snapshot_f12_0_a2_6, N_113_i_i_0, N_112_i_i_0, 
        start_snapshot_f12_0_a2_3, N_108_i_i_0, N_83_i_i_0, 
        N_111_i_i_0, N_82_i_i_0, \start_snapshot_f2_temp\, 
        counter_delta_snapshot_e12_i_0_o2_m6_e_6, 
        counter_delta_snapshot_e12_i_0_o2_m6_e_4, 
        counter_delta_snapshot_e12_i_0_o2_m6_e_5, 
        counter_delta_snapshot_e12_i_0_o2_m6_e_2, 
        un12_start_snapshot_fothers_temp_NE_5, 
        un12_start_snapshot_fothers_temp_NE_4, 
        un12_start_snapshot_fothers_temp_NE_11, 
        un12_start_snapshot_fothers_temp_NE_1, 
        un12_start_snapshot_fothers_temp_NE_0, 
        un12_start_snapshot_fothers_temp_NE_9, N_506_i, N_166_i_i, 
        un12_start_snapshot_fothers_temp_NE_7, N_133_i_i, 
        N_132_i_i, un12_start_snapshot_fothers_temp_NE_3, N_509_i, 
        N_164_i_i, N_510_i, N_135_i_i, 
        un12_start_snapshot_fothers_temp_NE_RNO_8, N_137_i_i, 
        counter_delta_f0_1_0_a2_12, counter_delta_f0_1_0_a2_1_0, 
        counter_delta_f0_1_0_a2_9, counter_delta_f0_1_0_a2_11, 
        counter_delta_f0_1_0_a2_6, counter_delta_f0_1_0_a2_5, 
        counter_delta_f0_1_0_a2_10, counter_delta_f0_1_0_a2_5_0, 
        counter_delta_f0_1_0_a2_0, N_272, 
        counter_delta_f0_1_0_a2_8_0, counter_delta_f0_1_0_a2_8_1, 
        counter_delta_f0_1_0_a2_3, counter_delta_f0_1_0_a2_2, 
        un1_start_snapshot_f22_i_a2_0_4, 
        un1_start_snapshot_f22_i_a2_0_3, 
        start_snapshot_f22_0_a2_11_0_a2_0, 
        \counter_delta_snapshot[17]_net_1\, start_snapshot_f12, 
        N_322, N_19, N_275, N_22_i_0, N_503, N_501, N_26, N_287, 
        N_288, N_6, N_486, N_488, N_8, N_480, N_482, 
        \counter_delta_snapshot_RNO[10]_net_1\, N_476, N_477, 
        \counter_delta_snapshot_RNO[9]_net_1\, N_471, N_472, 
        \counter_delta_snapshot_RNO[7]_net_1\, N_462, N_463, 
        \counter_delta_snapshot_RNO[6]_net_1\, N_457, N_458, 
        N_376_i_0, N_453, N_452, N_375_i_0, N_448, N_447, 
        \counter_delta_snapshot_RNO[3]_net_1\, N_442, N_443, N_54, 
        N_437, N_438, \counter_delta_snapshot_RNO[1]_net_1\, 
        N_433, counter_delta_snapshot_e1_i_0, N_435, N_263, N_259, 
        N_255, N_252, \counter_delta_snapshot_RNO[0]_net_1\, 
        N_505, counter_delta_snapshot_e24, N_192, N_193, N_194, 
        counter_delta_snapshot_e23, N_404, 
        counter_delta_snapshot_e22, N_186, N_187, N_188, 
        counter_delta_snapshot_e21, N_402, 
        \counter_delta_snapshot_RNO[20]_net_1\, N_180, N_181, 
        N_182, N_20, N_400, 
        \counter_delta_snapshot_RNO[17]_net_1\, N_171, N_172, 
        N_173, \counter_delta_snapshot_RNO[16]_net_1\, N_397, 
        N_390, N_504, N_383, \counter_delta_snapshot[1]_net_1\, 
        \counter_delta_snapshot[20]_net_1\, counter_delta_f0_1, 
        N_174, N_405, N_468, N_498, 
        \counter_delta_snapshot_RNO[18]_net_1\, N_175, N_176, 
        counter_delta_snapshot_e25, N_406, 
        \counter_delta_snapshot_RNO[8]_net_1\, N_467, 
        \counter_delta_snapshot_RNO[12]_net_1\, N_496, N_284, 
        counter_delta_snapshot_e26_0_0_0_tz, N_9, 
        counter_delta_snapshot_e26, N_425, N_21, N_23, N_107_i_i, 
        N_227, N_114_i_i, N_228, N_115_i_i, counter_delta_f0_n12, 
        counter_delta_f0_n13, counter_delta_f0_n14, 
        counter_delta_f0_n15, counter_delta_f0_n16, 
        counter_delta_f0_n17, counter_delta_f0_n18, N_11, 
        N_87_i_i, N_17, N_324_i, N_99_i_i, N_89_i_i, N_15, N_13, 
        N_117_i_i, N_116_i_i, N_230, N_229, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 


    \counter_delta_snapshot_RNO_1[11]\ : AOI1B
      port map(A => counter_delta_snapshot_e11_i_0_a2_0, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => N_294, Y
         => counter_delta_snapshot_e11_i_0_0);
    
    \counter_delta_snapshot_RNO[21]\ : OAI1
      port map(A => N_402, B => N_504_0, C => 
        counter_delta_snapshot_e21_0_0_0, Y => 
        counter_delta_snapshot_e21);
    
    \counter_delta_snapshot[19]\ : DFN1C0
      port map(D => N_20, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[19]_net_1\);
    
    start_snapshot_f0_RNO_1 : NOR3A
      port map(A => counter_delta_f0_1_0_a2_5_0, B => 
        counter_delta_f0_1_0_a2_0, C => N_272, Y => 
        counter_delta_f0_1_0_a2_10);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_6\ : NOR3C
      port map(A => N_133_i_i, B => N_132_i_i, C => 
        un12_start_snapshot_fothers_temp_NE_3, Y => 
        un12_start_snapshot_fothers_temp_NE_9);
    
    \counter_delta_f0_RNO[14]\ : AO1C
      port map(A => N_101, B => N_57_0, C => N_255, Y => 
        counter_delta_f0_n14);
    
    \op_eq.start_snapshot_f2_temp3_0_a2_RNO\ : OR2
      port map(A => start_snapshot_f22_11_i, B => 
        start_snapshot_f22_10, Y => 
        start_snapshot_f2_temp3_0_a2_0);
    
    \counter_delta_snapshot_RNO_0[17]\ : OR3C
      port map(A => N_397, B => 
        \counter_delta_snapshot[17]_net_1\, C => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_171);
    
    \counter_delta_snapshot_RNIP067[1]\ : NOR2
      port map(A => \counter_delta_snapshot[1]_net_1\, B => 
        \counter_delta_snapshot[0]_net_1\, Y => N_382);
    
    \counter_delta_f0_RNITCA8[6]\ : NOR2
      port map(A => \counter_delta_f0[7]_net_1\, B => 
        \counter_delta_f0[6]_net_1\, Y => 
        counter_delta_f0_1_0_a2_7);
    
    \counter_delta_snapshot_RNO_5[13]\ : OR2
      port map(A => \counter_delta_snapshot[13]_net_1\, B => 
        N_393, Y => counter_delta_snapshot_e13_i_0_a2_0);
    
    \counter_delta_snapshot_RNIKDF23[19]\ : OR3
      port map(A => N_398, B => 
        \counter_delta_snapshot[18]_net_1\, C => 
        \counter_delta_snapshot[19]_net_1\, Y => N_400);
    
    coarse_time_0_r_RNIGJTR4_0 : OR2B
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => un2_coarse_time_0, Y => N_504);
    
    \counter_delta_snapshot_RNIV4TS1[13]\ : NOR2A
      port map(A => N_393, B => 
        \counter_delta_snapshot[13]_net_1\, Y => N_394);
    
    \counter_delta_snapshot_RNO[19]\ : OAI1
      port map(A => N_400, B => N_504_0, C => 
        counter_delta_snapshot_e19_i_i_0, Y => N_20);
    
    \counter_delta_snapshot_RNO_1[2]\ : AO1A
      port map(A => counter_delta_snapshot_e2_i_a2_0, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => N_436, Y
         => counter_delta_snapshot_e2_i_0);
    
    \counter_delta_f0_RNO[11]\ : XA1A
      port map(A => N_67, B => \counter_delta_f0[11]_net_1\, C
         => N_57_0, Y => N_275);
    
    \counter_delta_f0_RNO_0[4]\ : AX1B
      port map(A => N_89, B => \counter_delta_f0[3]_net_1\, C => 
        \counter_delta_f0[4]_net_1\, Y => N_116_i_i);
    
    \counter_delta_f0_RNILJOA[20]\ : NOR3
      port map(A => \counter_delta_f0[14]_net_1\, B => 
        \counter_delta_f0[15]_net_1\, C => 
        \counter_delta_f0[20]_net_1\, Y => 
        counter_delta_f0_1_0_a2_3);
    
    \counter_delta_snapshot_RNO_1[12]\ : OR2
      port map(A => N_493, B => N_495, Y => 
        counter_delta_snapshot_e12_i_0_0);
    
    \counter_delta_snapshot_RNIIDER3[23]\ : OR3
      port map(A => N_402, B => 
        \counter_delta_snapshot[22]_net_1\, C => 
        \counter_delta_snapshot[23]_net_1\, Y => N_404);
    
    \counter_delta_f0_RNO[26]\ : XA1
      port map(A => N_80, B => \counter_delta_f0[26]_net_1\, C
         => N_57_0, Y => N_34);
    
    \counter_delta_snapshot_RNO_1[19]\ : OA1
      port map(A => N_398, B => 
        \counter_delta_snapshot[18]_net_1\, C => 
        \counter_delta_snapshot[19]_net_1\, Y => 
        counter_delta_snapshot_e19_i_i_a2_0);
    
    coarse_time_0_r_RNILJMD : NOR2A
      port map(A => coarse_time_0_c, B => \coarse_time_0_r\, Y
         => un2_coarse_time_0);
    
    \counter_delta_snapshot_RNO[5]\ : OR3C
      port map(A => N_453, B => counter_delta_snapshot_e5_i_0, C
         => N_452, Y => N_376_i_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_11\ : XNOR2
      port map(A => \counter_delta_snapshot[3]_net_1\, B => 
        delta_snapshot(3), Y => N_506_i);
    
    \counter_delta_snapshot[16]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[16]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[16]_net_1\);
    
    \counter_delta_snapshot_RNIRV6E4_0[23]\ : OR3B
      port map(A => \counter_delta_snapshot_e27_0_0_o2_m6_e_3\, B
         => counter_delta_snapshot_e27_0_0_o2_m6_e_2, C => N_398, 
        Y => counter_delta_snapshot_e27_0_0_o2_N_7_0);
    
    \counter_delta_snapshot_RNO_0[20]\ : OR3C
      port map(A => N_400, B => 
        \counter_delta_snapshot[20]_net_1\, C => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_180);
    
    \counter_delta_snapshot_RNIS3OS[7]\ : NOR2A
      port map(A => N_387, B => \counter_delta_snapshot[7]_net_1\, 
        Y => N_388);
    
    start_snapshot_f22_0_a2_RNO : OR2
      port map(A => start_snapshot_f22_0_a2_0, B => 
        start_snapshot_f22_11_i, Y => start_snapshot_f22_0_a2_1);
    
    \counter_delta_snapshot_RNO_1[16]\ : OR2B
      port map(A => counter_delta_snapshot_e16_i_i_a2_0, B => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_168);
    
    \counter_delta_snapshot_RNO_0[10]\ : NOR2
      port map(A => N_505, B => delta_snapshot(10), Y => N_476);
    
    \counter_delta_snapshot[25]\ : DFN1C0
      port map(D => counter_delta_snapshot_e25, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[25]_net_1\);
    
    \counter_delta_f0_RNO[7]\ : MX2
      port map(A => delta_f2_f0(7), B => N_89_i_i, S => N_57, Y
         => N_13);
    
    \counter_delta_snapshot_RNO_2[13]\ : NOR2A
      port map(A => counter_delta_snapshot_e13_i_0_a2_2_0, B => 
        N_504_0, Y => N_288);
    
    \counter_delta_snapshot_RNO_3[5]\ : OR2B
      port map(A => counter_delta_snapshot_e5_i_a2_0, B => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_450);
    
    counter_delta_snapshot_e12_i_0_a2 : NOR2A
      port map(A => counter_delta_snapshot_e27_0_0_o2_N_7_0, B
         => \counter_delta_snapshot_e12_i_0_a2_0\, Y => N_493);
    
    \counter_delta_snapshot[14]\ : DFN1C0
      port map(D => N_6, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[14]_net_1\);
    
    \counter_delta_snapshot_RNO_1[17]\ : OR2A
      port map(A => \counter_delta_snapshot[17]_net_1\, B => 
        un2_coarse_time_0, Y => N_172);
    
    \counter_delta_f0[14]\ : DFN1E0C0
      port map(D => counter_delta_f0_n14, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[14]_net_1\);
    
    \counter_delta_snapshot_RNO_0[2]\ : NOR2
      port map(A => N_505, B => delta_snapshot(2), Y => N_437);
    
    \counter_delta_f0_RNO[18]\ : AO1B
      port map(A => N_105, B => N_57, C => N_263, Y => 
        counter_delta_f0_n18);
    
    \counter_delta_snapshot_RNO[26]\ : AO1B
      port map(A => counter_delta_snapshot_e26_0_0_0_tz, B => 
        \counter_delta_snapshot[26]_net_1\, C => N_425, Y => 
        counter_delta_snapshot_e26);
    
    \counter_delta_snapshot_RNO[17]\ : OR3C
      port map(A => N_171, B => N_172, C => N_173, Y => 
        \counter_delta_snapshot_RNO[17]_net_1\);
    
    \counter_delta_snapshot[2]\ : DFN1C0
      port map(D => N_54, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[2]_net_1\);
    
    \counter_delta_f0_RNITVJ91[3]\ : NOR3A
      port map(A => counter_delta_f0lde_i_a2_0_1_2, B => N_89, C
         => \counter_delta_f0[3]_net_1\, Y => 
        counter_delta_f0lde_i_a2_0_1_3);
    
    \counter_delta_f0_RNIIVPK[4]\ : OR3
      port map(A => N_89, B => \counter_delta_f0[3]_net_1\, C => 
        \counter_delta_f0[4]_net_1\, Y => N_55);
    
    \counter_delta_snapshot_RNO_2[15]\ : NOR3B
      port map(A => N_395, B => 
        \counter_delta_snapshot[15]_net_1\, C => N_504_0, Y => 
        N_482);
    
    \counter_delta_snapshot_RNI5NLF2[16]\ : OR2
      port map(A => \counter_delta_snapshot[16]_net_1\, B => 
        N_396, Y => N_397);
    
    \counter_delta_f0_RNIU25H2[20]\ : OR2
      port map(A => \counter_delta_f0[20]_net_1\, B => N_106, Y
         => N_58);
    
    \counter_delta_snapshot_RNI71PA[2]\ : OR2A
      port map(A => N_382, B => \counter_delta_snapshot[2]_net_1\, 
        Y => N_383);
    
    \counter_delta_snapshot_RNO_2[14]\ : NOR3B
      port map(A => N_394, B => 
        \counter_delta_snapshot[14]_net_1\, C => N_504_0, Y => 
        N_488);
    
    \counter_delta_f0_RNO[20]\ : XA1A
      port map(A => \counter_delta_f0[20]_net_1\, B => N_106, C
         => N_57, Y => counter_delta_f0_n20);
    
    \counter_delta_snapshot_RNO_3[7]\ : NOR2A
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => counter_delta_snapshot_e7_i_a2_0, Y => N_460);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_5\ : NOR3C
      port map(A => N_506_i, B => N_166_i_i, C => 
        un12_start_snapshot_fothers_temp_NE_7, Y => 
        un12_start_snapshot_fothers_temp_NE_11);
    
    \counter_delta_snapshot[21]\ : DFN1C0
      port map(D => counter_delta_snapshot_e21, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[21]_net_1\);
    
    \counter_delta_f0_RNIPJ57[22]\ : OR2
      port map(A => \counter_delta_f0[23]_net_1\, B => 
        \counter_delta_f0[22]_net_1\, Y => 
        counter_delta_f0_1_0_a2_2);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_15\ : XNOR2
      port map(A => \counter_delta_snapshot[12]_net_1\, B => 
        delta_snapshot(12), Y => N_132_i_i);
    
    \counter_delta_f0[15]\ : DFN1E0C0
      port map(D => counter_delta_f0_n15, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[15]_net_1\);
    
    \counter_delta_snapshot_RNO_2[11]\ : OR2
      port map(A => N_505, B => delta_snapshot(11), Y => N_501);
    
    \counter_delta_f0_RNIBRBK1[12]\ : OR3
      port map(A => N_67, B => \counter_delta_f0[11]_net_1\, C
         => \counter_delta_f0[12]_net_1\, Y => N_99);
    
    \counter_delta_f0_RNI4JID2[19]\ : OR2A
      port map(A => N_105, B => \counter_delta_f0[19]_net_1\, Y
         => N_106);
    
    \counter_delta_snapshot_RNO[20]\ : OR3C
      port map(A => N_180, B => N_181, C => N_182, Y => 
        \counter_delta_snapshot_RNO[20]_net_1\);
    
    \counter_delta_snapshot_RNO_1[10]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[10]_net_1\, C => N_474, Y => 
        counter_delta_snapshot_e10_i_0);
    
    \counter_delta_snapshot_RNO[25]\ : OAI1
      port map(A => N_406, B => N_504, C => 
        counter_delta_snapshot_e25_0_0_0, Y => 
        counter_delta_snapshot_e25);
    
    \op_eq.start_snapshot_f2_temp3_0_a2\ : NOR2
      port map(A => un12_start_snapshot_fothers_temp_NE, B => 
        start_snapshot_f2_temp3_0_a2_0, Y => 
        start_snapshot_f2_temp3);
    
    \counter_delta_f0_RNIDC4T[6]\ : OR3
      port map(A => N_55, B => \counter_delta_f0[5]_net_1\, C => 
        \counter_delta_f0[6]_net_1\, Y => N_59);
    
    \counter_delta_f0_RNO_0[14]\ : OAI1
      port map(A => N_99, B => \counter_delta_f0[13]_net_1\, C
         => counter_delta_f0_n14_0_0_a2_0, Y => N_255);
    
    \counter_delta_snapshot_RNO[4]\ : NOR3C
      port map(A => N_448, B => counter_delta_snapshot_e4_i_0, C
         => N_447, Y => N_375_i_0);
    
    \counter_delta_snapshot[23]\ : DFN1C0
      port map(D => counter_delta_snapshot_e23, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[23]_net_1\);
    
    \counter_delta_snapshot_RNO_4[8]\ : NOR2
      port map(A => un2_coarse_time_0, B => 
        \counter_delta_snapshot[8]_net_1\, Y => N_466);
    
    \counter_delta_snapshot_RNO[23]\ : OAI1
      port map(A => N_404, B => N_504_0, C => 
        counter_delta_snapshot_e23_0_0_0, Y => 
        counter_delta_snapshot_e23);
    
    \counter_delta_snapshot[17]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[17]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[17]_net_1\);
    
    \counter_delta_f0[4]\ : DFN1E0C0
      port map(D => N_229, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[4]_net_1\);
    
    \counter_delta_f0_RNIVJ67[16]\ : NOR2
      port map(A => \counter_delta_f0[16]_net_1\, B => 
        \counter_delta_f0[17]_net_1\, Y => 
        counter_delta_f0_1_0_a2_8_0);
    
    counter_delta_snapshot_e27_0_0_o2_m6_e_3 : NOR2
      port map(A => \counter_delta_snapshot[23]_net_1\, B => 
        \counter_delta_snapshot[22]_net_1\, Y => 
        start_snapshot_f22_0_a2_11_0_a2_3_i);
    
    \counter_delta_f0[13]\ : DFN1E0C0
      port map(D => counter_delta_f0_n13, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[13]_net_1\);
    
    \counter_delta_snapshot_RNO_2[12]\ : NOR3A
      port map(A => \counter_delta_snapshot[12]_net_1\, B => 
        \counter_delta_snapshot_RNI0DDG1[7]_net_1\, C => N_504, Y
         => N_498);
    
    \counter_delta_f0_RNO_0[10]\ : AX1D
      port map(A => N_63, B => \counter_delta_f0[9]_net_1\, C => 
        \counter_delta_f0[10]_net_1\, Y => 
        counter_delta_f0_n10_0_i_0);
    
    \counter_delta_snapshot_RNO_2[19]\ : OR2A
      port map(A => \counter_delta_snapshot[19]_net_1\, B => 
        un2_coarse_time_0, Y => N_178);
    
    \counter_delta_f0_RNO_0[3]\ : XNOR2
      port map(A => \counter_delta_f0[3]_net_1\, B => N_89, Y => 
        N_115_i_i);
    
    \counter_delta_f0_RNI4NHR1[14]\ : OR3
      port map(A => N_99, B => \counter_delta_f0[13]_net_1\, C
         => \counter_delta_f0[14]_net_1\, Y => N_101);
    
    \counter_delta_snapshot_RNO_2[16]\ : NOR2B
      port map(A => \counter_delta_snapshot[16]_net_1\, B => 
        N_396, Y => counter_delta_snapshot_e16_i_i_a2_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_13\ : XA1A
      port map(A => delta_snapshot(6), B => 
        \counter_delta_snapshot[6]_net_1\, C => N_509_i, Y => 
        un12_start_snapshot_fothers_temp_NE_7);
    
    start_snapshot_fothers_temp : DFN1E0C0
      port map(D => N_7, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_284, Q => \start_snapshot_fothers_temp\);
    
    \counter_delta_snapshot_RNO_1[5]\ : OA1A
      port map(A => \counter_delta_snapshot_i[5]\, B => 
        un2_coarse_time_0_0, C => N_450, Y => 
        counter_delta_snapshot_e5_i_0);
    
    \counter_delta_snapshot_RNO_2[17]\ : OR2
      port map(A => N_504, B => N_398, Y => N_173);
    
    \counter_delta_snapshot_RNO[7]\ : NOR3
      port map(A => N_462, B => counter_delta_snapshot_e7_i_0, C
         => N_463, Y => \counter_delta_snapshot_RNO[7]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter_delta_snapshot[10]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[10]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[10]_net_1\);
    
    \counter_delta_f0_RNICPE51[8]\ : OR3
      port map(A => N_59, B => \counter_delta_f0[7]_net_1\, C => 
        \counter_delta_f0[8]_net_1\, Y => N_63);
    
    start_snapshot_f1_RNO_6 : XNOR2
      port map(A => \counter_delta_f0[4]_net_1\, B => 
        delta_f2_f1(4), Y => N_112_i_i_0);
    
    counter_delta_snapshot_e27_0_0_o2_m6_e_1_RNI4AT3 : AND2
      port map(A => start_snapshot_f22_0_a2_11_0_a2_3_i, B => 
        start_snapshot_f22_0_a2_11_0_a2_2_i, Y => 
        start_snapshot_f22_0_a2_11_0_a2_2_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_7\ : XNOR2
      port map(A => \counter_delta_snapshot[7]_net_1\, B => 
        delta_snapshot(7), Y => N_164_i_i);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \counter_delta_snapshot_RNO_0[6]\ : NOR2
      port map(A => N_505, B => delta_snapshot(6), Y => N_457);
    
    \counter_delta_f0_RNI3477[18]\ : NOR2
      port map(A => \counter_delta_f0[18]_net_1\, B => 
        \counter_delta_f0[19]_net_1\, Y => 
        counter_delta_f0_1_0_a2_8_1);
    
    \counter_delta_f0_RNI1DA8[8]\ : NOR2
      port map(A => \counter_delta_f0[8]_net_1\, B => 
        \counter_delta_f0[9]_net_1\, Y => 
        counter_delta_f0_1_0_a2_2_0);
    
    \counter_delta_snapshot[3]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[3]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[3]_net_1\);
    
    \counter_delta_f0_RNO_0[7]\ : XNOR2
      port map(A => \counter_delta_f0[7]_net_1\, B => N_59, Y => 
        N_89_i_i);
    
    \counter_delta_f0_RNIU767[26]\ : OR2
      port map(A => \counter_delta_f0[26]_net_1\, B => 
        \counter_delta_f0[24]_net_1\, Y => 
        counter_delta_f0_1_0_a2_0);
    
    \counter_delta_snapshot_RNI2DD92[15]\ : OR2A
      port map(A => N_395, B => 
        \counter_delta_snapshot[15]_net_1\, Y => N_396);
    
    \start_snapshot_f0\ : DFN1C0
      port map(D => counter_delta_f0_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => start_snapshot_f0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_3\ : XA1A
      port map(A => delta_snapshot(2), B => 
        \counter_delta_snapshot[2]_net_1\, C => N_510_i, Y => 
        un12_start_snapshot_fothers_temp_NE_4);
    
    \counter_delta_snapshot[12]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[12]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[12]_net_1\);
    
    start_snapshot_f0_RNO_0 : NOR3B
      port map(A => counter_delta_f0_1_0_a2_7, B => 
        counter_delta_f0_1_0_a2_6, C => counter_delta_f0_1_0_a2_5, 
        Y => counter_delta_f0_1_0_a2_11);
    
    \counter_delta_snapshot_RNO_0[0]\ : AXOI2
      port map(A => counter_delta_snapshot_e27_0_0_o2_N_7_0, B
         => un2_coarse_time_0_0, C => 
        \counter_delta_snapshot[0]_net_1\, Y => 
        counter_delta_snapshot_e0_i_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE\ : NAND2
      port map(A => un12_start_snapshot_fothers_temp_NE_12, B => 
        un12_start_snapshot_fothers_temp_NE_13, Y => 
        un12_start_snapshot_fothers_temp_NE);
    
    \counter_delta_snapshot_RNO_2[10]\ : NOR3A
      port map(A => \counter_delta_snapshot[10]_net_1\, B => 
        N_390, C => N_504_0, Y => N_477);
    
    \counter_delta_snapshot_RNI0DDG1[7]\ : OR3B
      port map(A => counter_delta_snapshot_e12_i_0_o2_m6_e_6, B
         => counter_delta_snapshot_e12_i_0_o2_m6_e_5, C => N_383, 
        Y => \counter_delta_snapshot_RNI0DDG1[7]_net_1\);
    
    \counter_delta_f0_RNO[25]\ : XA1A
      port map(A => N_66, B => \counter_delta_f0[25]_net_1\, C
         => N_57, Y => N_32);
    
    \counter_delta_snapshot_RNO[12]\ : NOR3
      port map(A => N_496, B => counter_delta_snapshot_e12_i_0_0, 
        C => N_498, Y => \counter_delta_snapshot_RNO[12]_net_1\);
    
    start_snapshot_f2_temp : DFN1C0
      port map(D => start_snapshot_f2_temp3, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \start_snapshot_f2_temp\);
    
    \counter_delta_f0[20]\ : DFN1E0C0
      port map(D => counter_delta_f0_n20, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[20]_net_1\);
    
    start_snapshot_f1_RNO_7 : XA1A
      port map(A => delta_f2_f1(2), B => 
        \counter_delta_f0[2]_net_1\, C => N_83_i_i_0, Y => 
        start_snapshot_f12_0_a2_3);
    
    \counter_delta_snapshot_RNO_4[13]\ : NOR2B
      port map(A => \counter_delta_snapshot[13]_net_1\, B => 
        N_393, Y => counter_delta_snapshot_e13_i_0_a2_2_0);
    
    \counter_delta_snapshot_RNO_0[1]\ : NOR2
      port map(A => N_505, B => delta_snapshot(1), Y => N_433);
    
    \counter_delta_f0[17]\ : DFN1E0C0
      port map(D => counter_delta_f0_n17, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[17]_net_1\);
    
    \counter_delta_f0_RNO_0[26]\ : NOR2
      port map(A => \counter_delta_f0[25]_net_1\, B => N_66, Y
         => N_80);
    
    \counter_delta_snapshot_RNO_4[15]\ : OR2
      port map(A => \counter_delta_snapshot[15]_net_1\, B => 
        N_395, Y => counter_delta_snapshot_e15_i_0_a2_0);
    
    counter_delta_snapshot_e12_i_0_a2_0 : NOR2
      port map(A => \counter_delta_snapshot[12]_net_1\, B => 
        un2_coarse_time_0_0, Y => N_495);
    
    \counter_delta_f0[2]\ : DFN1E0C0
      port map(D => N_227, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[2]_net_1\);
    
    \counter_delta_snapshot_RNO[18]\ : OR3C
      port map(A => N_174, B => N_175, C => N_176, Y => 
        \counter_delta_snapshot_RNO[18]_net_1\);
    
    \counter_delta_snapshot_RNINLU74[25]\ : OR2A
      port map(A => N_405, B => 
        \counter_delta_snapshot[25]_net_1\, Y => N_406);
    
    counter_delta_snapshot_e12_i_0_a2_RNO : OR2A
      port map(A => \counter_delta_snapshot_RNI0DDG1[7]_net_1\, B
         => \counter_delta_snapshot[12]_net_1\, Y => 
        \counter_delta_snapshot_e12_i_0_a2_0\);
    
    \counter_delta_f0_RNIJBBE[25]\ : NOR3
      port map(A => \counter_delta_f0[21]_net_1\, B => 
        \counter_delta_f0[25]_net_1\, C => 
        counter_delta_f0_1_0_a2_2, Y => 
        counter_delta_f0_1_0_a2_5_0);
    
    start_snapshot_f1_RNO_2 : XA1A
      port map(A => delta_f2_f1(1), B => 
        \counter_delta_f0[1]_net_1\, C => N_111_i_i_0, Y => 
        start_snapshot_f12_0_a2_1);
    
    \counter_delta_snapshot_RNO_4[14]\ : OR2
      port map(A => \counter_delta_snapshot[14]_net_1\, B => 
        N_394, Y => counter_delta_snapshot_e14_i_0_a2_0);
    
    \counter_delta_f0[21]\ : DFN1E0C0
      port map(D => N_276, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9_0, Q => \counter_delta_f0[21]_net_1\);
    
    \counter_delta_f0_RNO[1]\ : MX2
      port map(A => delta_f2_f0(1), B => N_107_i_i, S => N_57_0, 
        Y => N_23);
    
    \counter_delta_snapshot_RNI9IOI_0[26]\ : NOR3
      port map(A => \counter_delta_snapshot[25]_net_1\, B => 
        \counter_delta_snapshot[26]_net_1\, C => 
        \counter_delta_snapshot[24]_net_1\, Y => 
        \counter_delta_snapshot_e27_0_0_o2_m6_e_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \counter_delta_snapshot_RNO_1[9]\ : AO1A
      port map(A => counter_delta_snapshot_e9_i_a2_0, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => N_470, Y
         => counter_delta_snapshot_e9_i_0);
    
    \counter_delta_snapshot_RNO_4[2]\ : NOR2
      port map(A => un2_coarse_time_0, B => 
        \counter_delta_snapshot[2]_net_1\, Y => N_436);
    
    start_snapshot_f0_RNO_4 : NOR2A
      port map(A => \counter_delta_f0[0]_net_1\, B => 
        \counter_delta_f0[3]_net_1\, Y => 
        counter_delta_f0_1_0_a2_1_0);
    
    \counter_delta_snapshot_RNO_1[3]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[3]_net_1\, C => N_440, Y => 
        counter_delta_snapshot_e3_i_0);
    
    \counter_delta_snapshot_RNO_0[3]\ : NOR2
      port map(A => N_505, B => delta_snapshot(3), Y => N_442);
    
    \counter_delta_snapshot_RNI7OGC[16]\ : NOR2
      port map(A => \counter_delta_snapshot[16]_net_1\, B => 
        \counter_delta_snapshot[17]_net_1\, Y => 
        start_snapshot_f22_0_a2_11_0_a2_0);
    
    \counter_delta_snapshot_RNO_4[11]\ : OR2A
      port map(A => \counter_delta_snapshot_i[11]\, B => 
        un2_coarse_time_0, Y => N_294);
    
    \counter_delta_snapshot_RNO_1[23]\ : OAI1
      port map(A => N_402, B => 
        \counter_delta_snapshot[22]_net_1\, C => 
        counter_delta_snapshot_e23_0_0_a2_0, Y => N_189);
    
    \counter_delta_f0_RNIMF6D1[10]\ : OR3
      port map(A => N_63, B => \counter_delta_f0[9]_net_1\, C => 
        \counter_delta_f0[10]_net_1\, Y => N_67);
    
    \counter_delta_snapshot_RNIKFM14[24]\ : NOR2
      port map(A => \counter_delta_snapshot[24]_net_1\, B => 
        N_404, Y => N_405);
    
    \counter_delta_f0_RNO[16]\ : AO1C
      port map(A => N_103, B => N_57, C => N_259, Y => 
        counter_delta_f0_n16);
    
    \counter_delta_f0_RNIRALB3[3]\ : AO1B
      port map(A => counter_delta_f0lde_i_a2_0_1_3, B => N_322, C
         => sample_f0_val_0, Y => N_9_tz);
    
    \counter_delta_f0_RNO[8]\ : MX2
      port map(A => delta_f2_f0(8), B => N_99_i_i, S => N_57, Y
         => N_15);
    
    \counter_delta_snapshot_RNO_1[25]\ : OR2
      port map(A => counter_delta_snapshot_e25_0_0_a2_0, B => 
        N_405, Y => N_421);
    
    start_snapshot_f1_RNO_8 : XNOR2
      port map(A => \counter_delta_f0[3]_net_1\, B => 
        delta_f2_f1(3), Y => N_111_i_i_0);
    
    \counter_delta_snapshot_RNO[2]\ : NOR3
      port map(A => N_437, B => counter_delta_snapshot_e2_i_0, C
         => N_438, Y => N_54);
    
    \counter_delta_snapshot[26]\ : DFN1C0
      port map(D => counter_delta_snapshot_e26, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[26]_net_1\);
    
    \start_snapshot_f1\ : DFN1C0
      port map(D => start_snapshot_f12, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => start_snapshot_f1);
    
    \counter_delta_snapshot_RNIM1CE[3]\ : OR2
      port map(A => \counter_delta_snapshot[3]_net_1\, B => N_383, 
        Y => N_384);
    
    \counter_delta_snapshot_RNO_1[7]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[7]_net_1\, C => N_460, Y => 
        counter_delta_snapshot_e7_i_0);
    
    \counter_delta_snapshot_RNIV6LM1[12]\ : NOR2
      port map(A => \counter_delta_snapshot_RNI0DDG1[7]_net_1\, B
         => \counter_delta_snapshot[12]_net_1\, Y => N_393);
    
    \counter_delta_f0_RNO[5]\ : MX2
      port map(A => delta_f2_f0(5), B => N_117_i_i, S => N_57, Y
         => N_230);
    
    \counter_delta_snapshot_RNO_1[24]\ : OR2A
      port map(A => \counter_delta_snapshot[24]_net_1\, B => 
        un2_coarse_time_0, Y => N_193);
    
    \counter_delta_snapshot_RNO[6]\ : NOR3
      port map(A => N_457, B => counter_delta_snapshot_e6_i_0, C
         => N_458, Y => \counter_delta_snapshot_RNO[6]_net_1\);
    
    \counter_delta_snapshot[24]\ : DFN1C0
      port map(D => counter_delta_snapshot_e24, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[24]_net_1\);
    
    \counter_delta_snapshot_RNO_3[13]\ : NOR2A
      port map(A => counter_delta_snapshot_e27_0_0_o2_N_7_0, B
         => counter_delta_snapshot_e13_i_0_a2_0, Y => N_285);
    
    \counter_delta_f0_RNO[4]\ : MX2
      port map(A => delta_f2_f0(4), B => N_116_i_i, S => N_57, Y
         => N_229);
    
    \counter_delta_snapshot_RNO_3[3]\ : NOR3B
      port map(A => N_383, B => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, C => 
        \counter_delta_snapshot[3]_net_1\, Y => N_440);
    
    \counter_delta_snapshot_RNI55U31[9]\ : OR2A
      port map(A => N_389, B => \counter_delta_snapshot[9]_net_1\, 
        Y => N_390);
    
    \counter_delta_snapshot_RNO_1[21]\ : OAI1
      port map(A => N_400, B => 
        \counter_delta_snapshot[20]_net_1\, C => 
        counter_delta_snapshot_e21_0_0_a2_0, Y => N_183);
    
    start_snapshot_f1_RNO_9 : XNOR2
      port map(A => \counter_delta_f0[7]_net_1\, B => 
        delta_f2_f1(7), Y => N_82_i_i_0);
    
    \counter_delta_snapshot_RNIG4B01[8]\ : NOR2A
      port map(A => N_388, B => \counter_delta_snapshot[8]_net_1\, 
        Y => N_389);
    
    \counter_delta_f0[12]\ : DFN1E0C0
      port map(D => counter_delta_f0_n12, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[12]_net_1\);
    
    \counter_delta_f0_RNO_1[16]\ : NOR2B
      port map(A => \counter_delta_f0[16]_net_1\, B => N_57_0, Y
         => counter_delta_f0_n16_0_0_a2_0);
    
    \counter_delta_snapshot_RNO_3[15]\ : NOR2A
      port map(A => counter_delta_snapshot_e27_0_0_o2_N_7_0, B
         => counter_delta_snapshot_e15_i_0_a2_0, Y => N_478);
    
    \counter_delta_snapshot_RNO_1[6]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[6]_net_1\, C => N_455, Y => 
        counter_delta_snapshot_e6_i_0);
    
    \counter_delta_f0_RNO[10]\ : NOR2A
      port map(A => N_57_0, B => counter_delta_f0_n10_0_i_0, Y
         => N_19);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_12\ : XNOR2
      port map(A => \counter_delta_snapshot[9]_net_1\, B => 
        delta_snapshot(9), Y => N_166_i_i);
    
    \counter_delta_snapshot_RNO_2[8]\ : NOR3B
      port map(A => N_388, B => \counter_delta_snapshot[8]_net_1\, 
        C => N_504, Y => N_468);
    
    \counter_delta_f0_RNILRIL[10]\ : NOR3B
      port map(A => counter_delta_f0_1_0_a2_8_0, B => 
        counter_delta_f0_1_0_a2_8_1, C => 
        counter_delta_f0_1_0_a2_5, Y => 
        un1_start_snapshot_f22_i_a2_0_3);
    
    \counter_delta_snapshot_RNO_3[14]\ : NOR2A
      port map(A => counter_delta_snapshot_e27_0_0_o2_N_7_0, B
         => counter_delta_snapshot_e14_i_0_a2_0, Y => N_484);
    
    counter_delta_snapshot_e26_0_0_a2_1 : VCC
      port map(Y => N_425);
    
    \counter_delta_f0[3]\ : DFN1E0C0
      port map(D => N_228, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[3]_net_1\);
    
    \counter_delta_snapshot_RNO_0[8]\ : NOR2
      port map(A => N_505, B => delta_snapshot(8), Y => N_467);
    
    \counter_delta_f0_RNI2VU92[18]\ : NOR3
      port map(A => N_103, B => \counter_delta_f0[17]_net_1\, C
         => \counter_delta_f0[18]_net_1\, Y => N_105);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_10\ : XNOR2
      port map(A => \counter_delta_snapshot[1]_net_1\, B => 
        delta_snapshot(1), Y => N_137_i_i);
    
    \counter_delta_snapshot_RNO_0[4]\ : OR3A
      port map(A => \counter_delta_snapshot[4]_net_1\, B => N_384, 
        C => N_504, Y => N_448);
    
    \counter_delta_f0_RNO_0[8]\ : AX1B
      port map(A => N_59, B => \counter_delta_f0[7]_net_1\, C => 
        \counter_delta_f0[8]_net_1\, Y => N_99_i_i);
    
    \counter_delta_f0[24]\ : DFN1E0C0
      port map(D => N_30, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[24]_net_1\);
    
    \counter_delta_snapshot_RNO_1[22]\ : OR2A
      port map(A => \counter_delta_snapshot[22]_net_1\, B => 
        un2_coarse_time_0, Y => N_187);
    
    \counter_delta_f0_RNO[23]\ : XA1A
      port map(A => N_62, B => \counter_delta_f0[23]_net_1\, C
         => N_57, Y => N_28);
    
    \counter_delta_snapshot_RNO_3[11]\ : NOR2B
      port map(A => \counter_delta_snapshot_i[11]\, B => N_391, Y
         => counter_delta_snapshot_e11_i_0_a2_0);
    
    \counter_delta_snapshot_RNO_2[1]\ : NOR3A
      port map(A => \counter_delta_snapshot[1]_net_1\, B => 
        \counter_delta_snapshot[0]_net_1\, C => N_504, Y => N_435);
    
    \counter_delta_f0_RNO_0[6]\ : AX1B
      port map(A => N_55, B => \counter_delta_f0[5]_net_1\, C => 
        \counter_delta_f0[6]_net_1\, Y => N_87_i_i);
    
    \counter_delta_f0_RNIAF4P[20]\ : NOR3A
      port map(A => counter_delta_f0_1_0_a2_3, B => 
        counter_delta_f0_1_0_a2_0, C => N_272, Y => 
        un1_start_snapshot_f22_i_a2_0_4);
    
    start_snapshot_f0_RNO_5 : NOR3C
      port map(A => counter_delta_f0_1_0_a2_8_0, B => 
        counter_delta_f0_1_0_a2_8_1, C => 
        counter_delta_f0_1_0_a2_3, Y => counter_delta_f0_1_0_a2_9);
    
    \counter_delta_f0_RNO_0[2]\ : AX1B
      port map(A => \counter_delta_f0[0]_net_1\, B => 
        \counter_delta_f0[1]_net_1\, C => 
        \counter_delta_f0[2]_net_1\, Y => N_114_i_i);
    
    \counter_delta_snapshot_RNO[22]\ : OR3C
      port map(A => N_186, B => N_187, C => N_188, Y => 
        counter_delta_snapshot_e22);
    
    \counter_delta_snapshot_RNO[1]\ : NOR3
      port map(A => N_433, B => counter_delta_snapshot_e1_i_0, C
         => N_435, Y => \counter_delta_snapshot_RNO[1]_net_1\);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_4\ : XA1A
      port map(A => delta_snapshot(0), B => 
        \counter_delta_snapshot[0]_net_1\, C => N_137_i_i, Y => 
        un12_start_snapshot_fothers_temp_NE_0);
    
    \counter_delta_snapshot_RNO[14]\ : NOR3
      port map(A => N_486, B => counter_delta_snapshot_e14_i_0_0, 
        C => N_488, Y => N_6);
    
    start_snapshot_fothers_temp_RNI1HGO3 : NOR2B
      port map(A => N_57_0, B => N_9_tz, Y => N_9_0);
    
    \counter_delta_snapshot_RNO_2[7]\ : NOR3B
      port map(A => N_387, B => \counter_delta_snapshot[7]_net_1\, 
        C => N_504_0, Y => N_463);
    
    \counter_delta_f0_RNO[3]\ : MX2
      port map(A => delta_f2_f0(3), B => N_115_i_i, S => N_57_0, 
        Y => N_228);
    
    \counter_delta_snapshot_RNO_2[23]\ : NOR2B
      port map(A => \counter_delta_snapshot[23]_net_1\, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, Y => 
        counter_delta_snapshot_e23_0_0_a2_0);
    
    \start_snapshot_f2\ : DFN1C0
      port map(D => N_7, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        start_snapshot_f2);
    
    start_snapshot_fothers_temp_RNI66RC : OAI1
      port map(A => N_7, B => \start_snapshot_fothers_temp\, C
         => sample_f2_val, Y => N_57_0);
    
    \counter_delta_snapshot_RNO_2[6]\ : NOR3A
      port map(A => \counter_delta_snapshot[6]_net_1\, B => N_386, 
        C => N_504_0, Y => N_458);
    
    \counter_delta_f0_RNILEAO2[22]\ : OR3
      port map(A => N_58, B => \counter_delta_f0[21]_net_1\, C
         => \counter_delta_f0[22]_net_1\, Y => N_62);
    
    \counter_delta_f0[25]\ : DFN1E0C0
      port map(D => N_32, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[25]_net_1\);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_1\ : XA1
      port map(A => delta_snapshot(5), B => 
        \counter_delta_snapshot_i[5]\, C => N_164_i_i, Y => 
        un12_start_snapshot_fothers_temp_NE_5);
    
    \counter_delta_snapshot_RNIRV6E4[23]\ : OR3B
      port map(A => \counter_delta_snapshot_e27_0_0_o2_m6_e_3\, B
         => counter_delta_snapshot_e27_0_0_o2_m6_e_2, C => N_398, 
        Y => \counter_delta_snapshot_RNIRV6E4[23]_net_1\);
    
    \counter_delta_snapshot_RNO_2[25]\ : OR2B
      port map(A => \counter_delta_snapshot[25]_net_1\, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, Y => 
        counter_delta_snapshot_e25_0_0_a2_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_9\ : XNOR2
      port map(A => \counter_delta_snapshot[10]_net_1\, B => 
        delta_snapshot(10), Y => N_510_i);
    
    \counter_delta_f0_RNO[9]\ : MX2
      port map(A => delta_f2_f0(9), B => N_324_i, S => N_57, Y
         => N_17);
    
    \counter_delta_f0_RNINJ57[12]\ : OR2
      port map(A => \counter_delta_f0[13]_net_1\, B => 
        \counter_delta_f0[12]_net_1\, Y => N_272);
    
    \counter_delta_f0[16]\ : DFN1E0C0
      port map(D => counter_delta_f0_n16, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[16]_net_1\);
    
    \counter_delta_snapshot_RNO_2[24]\ : OR2A
      port map(A => N_405, B => N_504, Y => N_194);
    
    \counter_delta_snapshot_RNIT7FC[21]\ : OR2
      port map(A => \counter_delta_snapshot[21]_net_1\, B => 
        \counter_delta_snapshot[20]_net_1\, Y => 
        start_snapshot_f22_0_a2_11_0_a2_1);
    
    start_snapshot_f0_RNO_3 : NOR3A
      port map(A => N_273, B => \counter_delta_f0[2]_net_1\, C
         => \counter_delta_f0[1]_net_1\, Y => 
        counter_delta_f0_1_0_a2_6);
    
    \counter_delta_snapshot_RNO_3[8]\ : OR2
      port map(A => \counter_delta_snapshot[8]_net_1\, B => N_388, 
        Y => counter_delta_snapshot_e8_i_a2_0);
    
    \counter_delta_snapshot_RNIN2IL[5]\ : OR2A
      port map(A => \counter_delta_snapshot_i[5]\, B => N_385, Y
         => N_386);
    
    \counter_delta_snapshot_RNO_3[9]\ : OR2
      port map(A => \counter_delta_snapshot[9]_net_1\, B => N_389, 
        Y => counter_delta_snapshot_e9_i_a2_0);
    
    \counter_delta_snapshot_RNO_2[3]\ : NOR3A
      port map(A => \counter_delta_snapshot[3]_net_1\, B => N_383, 
        C => N_504, Y => N_443);
    
    \counter_delta_f0_RNO[19]\ : AO1C
      port map(A => N_106, B => N_57, C => N_265, Y => 
        counter_delta_f0_n19);
    
    start_snapshot_f1_RNO_11 : XNOR2
      port map(A => \counter_delta_f0[8]_net_1\, B => 
        delta_f2_f1(8), Y => N_83_i_i_0);
    
    \counter_delta_f0_RNO_0[1]\ : XNOR2
      port map(A => \counter_delta_f0[1]_net_1\, B => 
        \counter_delta_f0[0]_net_1\, Y => N_107_i_i);
    
    \counter_delta_f0_RNIRIFC[2]\ : OR3
      port map(A => \counter_delta_f0[0]_net_1\, B => 
        \counter_delta_f0[1]_net_1\, C => 
        \counter_delta_f0[2]_net_1\, Y => N_89);
    
    \counter_delta_snapshot_RNO_2[21]\ : NOR2B
      port map(A => \counter_delta_snapshot[21]_net_1\, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, Y => 
        counter_delta_snapshot_e21_0_0_a2_0);
    
    \counter_delta_snapshot[20]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[20]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[20]_net_1\);
    
    \counter_delta_f0_RNO_0[22]\ : AX1D
      port map(A => N_58, B => \counter_delta_f0[21]_net_1\, C
         => \counter_delta_f0[22]_net_1\, Y => N_86_i);
    
    \counter_delta_f0[0]\ : DFN1E0C0
      port map(D => N_21, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9_0, Q => \counter_delta_f0[0]_net_1\);
    
    \counter_delta_f0[23]\ : DFN1E0C0
      port map(D => N_28, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[23]_net_1\);
    
    \counter_delta_snapshot_RNI9KJK[7]\ : NOR3A
      port map(A => counter_delta_snapshot_e12_i_0_o2_m6_e_4, B
         => \counter_delta_snapshot[8]_net_1\, C => 
        \counter_delta_snapshot[7]_net_1\, Y => 
        counter_delta_snapshot_e12_i_0_o2_m6_e_6);
    
    \counter_delta_f0_RNO[22]\ : NOR2A
      port map(A => N_57, B => N_86_i, Y => N_277);
    
    \counter_delta_f0[8]\ : DFN1E0C0
      port map(D => N_15, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[8]_net_1\);
    
    \counter_delta_snapshot_RNO_1[20]\ : OR2A
      port map(A => \counter_delta_snapshot[20]_net_1\, B => 
        un2_coarse_time_0, Y => N_181);
    
    \counter_delta_snapshot_RNO_0[9]\ : NOR2
      port map(A => N_505, B => delta_snapshot(9), Y => N_471);
    
    \counter_delta_f0_RNO_1[18]\ : NOR2B
      port map(A => \counter_delta_f0[18]_net_1\, B => N_57_0, Y
         => counter_delta_f0_n18_0_0_a2_0);
    
    start_snapshot_f1_RNO : NOR3C
      port map(A => start_snapshot_f12_0_a2_7, B => 
        start_snapshot_f12_0_a2_6, C => N_322, Y => 
        start_snapshot_f12);
    
    \counter_delta_f0_RNO[2]\ : MX2
      port map(A => delta_f2_f0(2), B => N_114_i_i, S => N_57_0, 
        Y => N_227);
    
    start_snapshot_f0_RNO_2 : NOR3C
      port map(A => counter_delta_f0_1_0_a2_2_0, B => 
        counter_delta_f0_1_0_a2_1_0, C => 
        counter_delta_f0_1_0_a2_9, Y => 
        counter_delta_f0_1_0_a2_12);
    
    \counter_delta_snapshot_RNO_1[4]\ : OA1
      port map(A => \counter_delta_snapshot[4]_net_1\, B => 
        un2_coarse_time_0_0, C => N_445, Y => 
        counter_delta_snapshot_e4_i_0);
    
    \counter_delta_snapshot_RNIGN0H[11]\ : NOR3B
      port map(A => \counter_delta_snapshot_i[11]\, B => 
        counter_delta_snapshot_e12_i_0_o2_m6_e_2, C => 
        \counter_delta_snapshot[3]_net_1\, Y => 
        counter_delta_snapshot_e12_i_0_o2_m6_e_5);
    
    \counter_delta_snapshot_RNIAA8V[23]\ : NOR3A
      port map(A => \counter_delta_snapshot_e27_0_0_o2_m6_e_1\, B
         => \counter_delta_snapshot[22]_net_1\, C => 
        \counter_delta_snapshot[23]_net_1\, Y => 
        \counter_delta_snapshot_e27_0_0_o2_m6_e_3\);
    
    coarse_time_0_r_RNIGJTR4 : OR2B
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => un2_coarse_time_0_0, Y => N_504_0);
    
    start_snapshot_f0_RNO : NOR3C
      port map(A => counter_delta_f0_1_0_a2_11, B => 
        counter_delta_f0_1_0_a2_10, C => 
        counter_delta_f0_1_0_a2_12, Y => counter_delta_f0_1);
    
    \counter_delta_snapshot_RNO_2[22]\ : OR3
      port map(A => N_402, B => 
        \counter_delta_snapshot[22]_net_1\, C => N_504, Y => 
        N_188);
    
    \counter_delta_snapshot_RNO[9]\ : NOR3
      port map(A => N_471, B => counter_delta_snapshot_e9_i_0, C
         => N_472, Y => \counter_delta_snapshot_RNO[9]_net_1\);
    
    start_snapshot_f1_RNO_5 : XNOR2
      port map(A => \counter_delta_f0[5]_net_1\, B => 
        delta_f2_f1(5), Y => N_113_i_i_0);
    
    \counter_delta_f0[1]\ : DFN1E0C0
      port map(D => N_23, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9_0, Q => \counter_delta_f0[1]_net_1\);
    
    \counter_delta_snapshot_RNI95UL2[17]\ : OR2
      port map(A => \counter_delta_snapshot[17]_net_1\, B => 
        N_397, Y => N_398);
    
    \counter_delta_snapshot[22]\ : DFN1C0
      port map(D => counter_delta_snapshot_e22, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \counter_delta_snapshot[22]_net_1\);
    
    \counter_delta_f0_RNO[15]\ : XA1A
      port map(A => \counter_delta_f0[15]_net_1\, B => N_101, C
         => N_57_0, Y => counter_delta_f0_n15);
    
    \counter_delta_f0[19]\ : DFN1E0C0
      port map(D => counter_delta_f0_n19, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[19]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \counter_delta_snapshot_RNO_0[5]\ : OR3
      port map(A => N_385, B => \counter_delta_snapshot_i[5]\, C
         => N_504_0, Y => N_453);
    
    \counter_delta_f0_RNO[24]\ : NOR2A
      port map(A => N_57, B => N_98_i, Y => N_30);
    
    \counter_delta_snapshot_RNO[3]\ : NOR3
      port map(A => N_442, B => counter_delta_snapshot_e3_i_0, C
         => N_443, Y => \counter_delta_snapshot_RNO[3]_net_1\);
    
    \counter_delta_f0_RNO_0[16]\ : OAI1
      port map(A => N_101, B => \counter_delta_f0[15]_net_1\, C
         => counter_delta_f0_n16_0_0_a2_0, Y => N_259);
    
    \counter_delta_snapshot[6]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[6]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[6]_net_1\);
    
    \counter_delta_f0[18]\ : DFN1E0C0
      port map(D => counter_delta_f0_n18, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_9_0, Q => \counter_delta_f0[18]_net_1\);
    
    \counter_delta_snapshot_RNO_3[10]\ : NOR3B
      port map(A => N_390, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => 
        \counter_delta_snapshot[10]_net_1\, Y => N_474);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_8\ : XOR2
      port map(A => \counter_delta_snapshot_i[11]\, B => 
        delta_snapshot(11), Y => 
        un12_start_snapshot_fothers_temp_NE_RNO_8);
    
    start_snapshot_fothers_temp_RNI66RC_0 : OAI1
      port map(A => N_7, B => \start_snapshot_fothers_temp\, C
         => sample_f2_val, Y => N_57);
    
    \counter_delta_f0[6]\ : DFN1E0C0
      port map(D => N_11, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[6]_net_1\);
    
    \counter_delta_snapshot[8]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[8]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[8]_net_1\);
    
    \counter_delta_snapshot_RNO_0[18]\ : OR3C
      port map(A => N_398, B => 
        \counter_delta_snapshot[18]_net_1\, C => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_174);
    
    counter_delta_snapshot_e27_0_0_o2_m6_e_1_RNI8ATS : OR3B
      port map(A => start_snapshot_f22_0_a2_11_0_a2_0, B => 
        start_snapshot_f22_0_a2_11_0_a2_2_0, C => 
        start_snapshot_f22_0_a2_11_0_a2_1, Y => 
        start_snapshot_f22_11_i);
    
    \counter_delta_snapshot_RNI2JDD[4]\ : NOR3
      port map(A => \counter_delta_snapshot[10]_net_1\, B => 
        \counter_delta_snapshot[4]_net_1\, C => 
        \counter_delta_snapshot[9]_net_1\, Y => 
        counter_delta_snapshot_e12_i_0_o2_m6_e_4);
    
    start_snapshot_f1_RNO_0 : NOR3C
      port map(A => start_snapshot_f12_0_a2_1, B => 
        start_snapshot_f12_0_a2_0, C => start_snapshot_f12_0_a2_4, 
        Y => start_snapshot_f12_0_a2_7);
    
    \counter_delta_f0_RNO[21]\ : XA1A
      port map(A => N_58, B => \counter_delta_f0[21]_net_1\, C
         => N_57, Y => N_276);
    
    \counter_delta_snapshot_RNO_4[7]\ : OR2
      port map(A => \counter_delta_snapshot[7]_net_1\, B => N_387, 
        Y => counter_delta_snapshot_e7_i_a2_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_17\ : XNOR2
      port map(A => \counter_delta_snapshot[8]_net_1\, B => 
        delta_snapshot(8), Y => N_509_i);
    
    \counter_delta_f0_RNIIM2T1[25]\ : NOR3C
      port map(A => un1_start_snapshot_f22_i_a2_0_3, B => 
        counter_delta_f0_1_0_a2_5_0, C => 
        un1_start_snapshot_f22_i_a2_0_4, Y => N_322);
    
    \counter_delta_snapshot[4]\ : DFN1C0
      port map(D => N_375_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => \counter_delta_snapshot[4]_net_1\);
    
    \counter_delta_snapshot_RNI935P[6]\ : NOR2
      port map(A => \counter_delta_snapshot[6]_net_1\, B => N_386, 
        Y => N_387);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_0\ : NOR3C
      port map(A => un12_start_snapshot_fothers_temp_NE_5, B => 
        un12_start_snapshot_fothers_temp_NE_4, C => 
        un12_start_snapshot_fothers_temp_NE_11, Y => 
        un12_start_snapshot_fothers_temp_NE_13);
    
    \counter_delta_snapshot_RNO[24]\ : OR3C
      port map(A => N_192, B => N_193, C => N_194, Y => 
        counter_delta_snapshot_e24);
    
    \counter_delta_f0_RNO_1[12]\ : NOR2B
      port map(A => \counter_delta_f0[12]_net_1\, B => N_57_0, Y
         => counter_delta_f0_n12_0_0_a2_0);
    
    \counter_delta_f0_RNIJ357[10]\ : OR2
      port map(A => \counter_delta_f0[11]_net_1\, B => 
        \counter_delta_f0[10]_net_1\, Y => 
        counter_delta_f0_1_0_a2_5);
    
    \counter_delta_snapshot[15]\ : DFN1C0
      port map(D => N_8, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[15]_net_1\);
    
    \counter_delta_snapshot_RNO_1[1]\ : OA1C
      port map(A => un2_coarse_time_0, B => 
        \counter_delta_snapshot[0]_net_1\, C => 
        \counter_delta_snapshot[1]_net_1\, Y => 
        counter_delta_snapshot_e1_i_0);
    
    \counter_delta_snapshot_RNO_3[2]\ : OR2
      port map(A => \counter_delta_snapshot[2]_net_1\, B => N_382, 
        Y => counter_delta_snapshot_e2_i_a2_0);
    
    start_snapshot_fothers_temp_RNI1HGO3_0 : NOR2B
      port map(A => N_57_0, B => N_9_tz, Y => N_9);
    
    \counter_delta_f0[9]\ : DFN1E0C0
      port map(D => N_17, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[9]_net_1\);
    
    \counter_delta_snapshot_RNO[0]\ : OA1B
      port map(A => delta_snapshot(0), B => N_505, C => 
        counter_delta_snapshot_e0_i_0, Y => 
        \counter_delta_snapshot_RNO[0]_net_1\);
    
    start_snapshot_f1_RNO_10 : XNOR2
      port map(A => \counter_delta_f0[0]_net_1\, B => 
        delta_f2_f1(0), Y => N_108_i_i_0);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO\ : NOR3C
      port map(A => un12_start_snapshot_fothers_temp_NE_1, B => 
        un12_start_snapshot_fothers_temp_NE_0, C => 
        un12_start_snapshot_fothers_temp_NE_9, Y => 
        un12_start_snapshot_fothers_temp_NE_12);
    
    \counter_delta_snapshot_RNO_2[20]\ : OR3
      port map(A => N_400, B => 
        \counter_delta_snapshot[20]_net_1\, C => N_504, Y => 
        N_182);
    
    \counter_delta_snapshot_RNO_4[5]\ : NOR2B
      port map(A => \counter_delta_snapshot_i[5]\, B => N_385, Y
         => counter_delta_snapshot_e5_i_a2_0);
    
    \counter_delta_snapshot_RNO_1[18]\ : OR2A
      port map(A => \counter_delta_snapshot[18]_net_1\, B => 
        un2_coarse_time_0, Y => N_175);
    
    \counter_delta_f0_RNO_0[9]\ : XNOR2
      port map(A => \counter_delta_f0[9]_net_1\, B => N_63, Y => 
        N_324_i);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_2\ : XA1A
      port map(A => delta_snapshot(4), B => 
        \counter_delta_snapshot[4]_net_1\, C => 
        un12_start_snapshot_fothers_temp_NE_RNO_8, Y => 
        un12_start_snapshot_fothers_temp_NE_1);
    
    \counter_delta_snapshot_RNI62VH[4]\ : OR2
      port map(A => \counter_delta_snapshot[4]_net_1\, B => N_384, 
        Y => N_385);
    
    \counter_delta_snapshot[11]\ : DFN1P0
      port map(D => N_22_i_0, CLK => HCLK_c, PRE => HRESETn_c, Q
         => \counter_delta_snapshot_i[11]\);
    
    \counter_delta_snapshot_RNO_4[9]\ : NOR2
      port map(A => un2_coarse_time_0, B => 
        \counter_delta_snapshot[9]_net_1\, Y => N_470);
    
    \counter_delta_f0_RNO_0[5]\ : XNOR2
      port map(A => \counter_delta_f0[5]_net_1\, B => N_55, Y => 
        N_117_i_i);
    
    \counter_delta_snapshot_RNI07532[14]\ : NOR2A
      port map(A => N_394, B => 
        \counter_delta_snapshot[14]_net_1\, Y => N_395);
    
    \counter_delta_snapshot_RNO_1[8]\ : AO1A
      port map(A => counter_delta_snapshot_e8_i_a2_0, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => N_466, Y
         => counter_delta_snapshot_e8_i_0);
    
    \counter_delta_snapshot_RNO_2[5]\ : OR2
      port map(A => N_505, B => delta_snapshot(5), Y => N_452);
    
    \counter_delta_snapshot_RNO[11]\ : OR3C
      port map(A => N_503, B => counter_delta_snapshot_e11_i_0_0, 
        C => N_501, Y => N_22_i_0);
    
    \counter_delta_snapshot[18]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[18]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[18]_net_1\);
    
    \counter_delta_f0_RNO_0[19]\ : OR3B
      port map(A => N_57_0, B => \counter_delta_f0[19]_net_1\, C
         => N_105, Y => N_265);
    
    \counter_delta_f0_RNO_0[18]\ : OAI1
      port map(A => N_103, B => \counter_delta_f0[17]_net_1\, C
         => counter_delta_f0_n18_0_0_a2_0, Y => N_263);
    
    \counter_delta_snapshot_RNO_2[2]\ : NOR3B
      port map(A => N_382, B => \counter_delta_snapshot[2]_net_1\, 
        C => N_504, Y => N_438);
    
    \counter_delta_snapshot[13]\ : DFN1C0
      port map(D => N_26, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[13]_net_1\);
    
    \counter_delta_snapshot_RNO_2[4]\ : OR2
      port map(A => N_505, B => delta_snapshot(4), Y => N_447);
    
    \counter_delta_snapshot_RNI9IOI[26]\ : OR3
      port map(A => \counter_delta_snapshot[25]_net_1\, B => 
        \counter_delta_snapshot[26]_net_1\, C => 
        \counter_delta_snapshot[24]_net_1\, Y => 
        start_snapshot_f22_10);
    
    \counter_delta_snapshot_RNI2N5A1[10]\ : OR2
      port map(A => \counter_delta_snapshot[10]_net_1\, B => 
        N_390, Y => N_391);
    
    \counter_delta_f0_RNO[17]\ : XA1A
      port map(A => \counter_delta_f0[17]_net_1\, B => N_103, C
         => N_57, Y => counter_delta_f0_n17);
    
    \counter_delta_snapshot_RNI3167[5]\ : NOR2A
      port map(A => \counter_delta_snapshot_i[5]\, B => 
        \counter_delta_snapshot[6]_net_1\, Y => 
        counter_delta_snapshot_e12_i_0_o2_m6_e_2);
    
    \counter_delta_snapshot_RNO_0[23]\ : OA1A
      port map(A => \counter_delta_snapshot[23]_net_1\, B => 
        un2_coarse_time_0_0, C => N_189, Y => 
        counter_delta_snapshot_e23_0_0_0);
    
    \counter_delta_f0_RNO[13]\ : XA1A
      port map(A => \counter_delta_f0[13]_net_1\, B => N_99, C
         => N_57_0, Y => counter_delta_f0_n13);
    
    \counter_delta_snapshot_RNO_0[13]\ : NOR2
      port map(A => N_505, B => delta_snapshot(13), Y => N_287);
    
    \counter_delta_snapshot_RNO[8]\ : NOR3
      port map(A => N_467, B => counter_delta_snapshot_e8_i_0, C
         => N_468, Y => \counter_delta_snapshot_RNO[8]_net_1\);
    
    \counter_delta_f0_RNO_0[24]\ : AX1D
      port map(A => N_62, B => \counter_delta_f0[23]_net_1\, C
         => \counter_delta_f0[24]_net_1\, Y => N_98_i);
    
    coarse_time_0_r_RNILJMD_0 : NOR2A
      port map(A => coarse_time_0_c, B => \coarse_time_0_r\, Y
         => un2_coarse_time_0_0);
    
    start_snapshot_f22_0_a2_RNO_0 : OR2
      port map(A => \start_snapshot_f2_temp\, B => 
        start_snapshot_f22_10, Y => start_snapshot_f22_0_a2_0);
    
    \counter_delta_f0_RNO[0]\ : MX2B
      port map(A => delta_f2_f0(0), B => 
        \counter_delta_f0[0]_net_1\, S => N_57_0, Y => N_21);
    
    coarse_time_0_r_RNIGJTR4_1 : OR2A
      port map(A => un2_coarse_time_0, B => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_505);
    
    \counter_delta_snapshot[1]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[1]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[1]_net_1\);
    
    \counter_delta_f0[22]\ : DFN1E0C0
      port map(D => N_277, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[22]_net_1\);
    
    \counter_delta_snapshot_RNO_0[25]\ : OA1A
      port map(A => \counter_delta_snapshot[25]_net_1\, B => 
        un2_coarse_time_0_0, C => N_421, Y => 
        counter_delta_snapshot_e25_0_0_0);
    
    \counter_delta_f0_RNI13O22[16]\ : OR3
      port map(A => N_101, B => \counter_delta_f0[15]_net_1\, C
         => \counter_delta_f0[16]_net_1\, Y => N_103);
    
    \counter_delta_snapshot_RNO_0[15]\ : NOR2
      port map(A => N_505, B => delta_snapshot(15), Y => N_480);
    
    \counter_delta_snapshot_RNO_0[24]\ : OR3C
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => \counter_delta_snapshot[24]_net_1\, C => N_404, Y
         => N_192);
    
    \counter_delta_snapshot_RNO_0[14]\ : NOR2
      port map(A => N_505, B => delta_snapshot(14), Y => N_486);
    
    start_snapshot_fothers_temp_RNO : NOR3B
      port map(A => N_322, B => counter_delta_f0lde_i_a2_0_1_3, C
         => N_7, Y => N_284);
    
    \counter_delta_snapshot_RNIHLUE3[21]\ : OR3
      port map(A => N_400, B => 
        \counter_delta_snapshot[20]_net_1\, C => 
        \counter_delta_snapshot[21]_net_1\, Y => N_402);
    
    \counter_delta_snapshot_RNI8G0P[19]\ : NOR3
      port map(A => \counter_delta_snapshot[18]_net_1\, B => 
        \counter_delta_snapshot[19]_net_1\, C => 
        start_snapshot_f22_0_a2_11_0_a2_1, Y => 
        counter_delta_snapshot_e27_0_0_o2_m6_e_2);
    
    \counter_delta_snapshot_RNO[16]\ : OAI1
      port map(A => N_397, B => N_504_0, C => 
        counter_delta_snapshot_e16_i_i_0, Y => 
        \counter_delta_snapshot_RNO[16]_net_1\);
    
    \counter_delta_f0_RNIN6VO[4]\ : NOR3C
      port map(A => counter_delta_f0_1_0_a2_7, B => N_273, C => 
        counter_delta_f0_1_0_a2_2_0, Y => 
        counter_delta_f0lde_i_a2_0_1_2);
    
    \counter_delta_f0[7]\ : DFN1E0C0
      port map(D => N_13, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[7]_net_1\);
    
    \counter_delta_snapshot_RNO_0[21]\ : OA1A
      port map(A => \counter_delta_snapshot[21]_net_1\, B => 
        un2_coarse_time_0, C => N_183, Y => 
        counter_delta_snapshot_e21_0_0_0);
    
    \counter_delta_f0[5]\ : DFN1E0C0
      port map(D => N_230, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[5]_net_1\);
    
    coarse_time_0_r : DFN1C0
      port map(D => coarse_time_0_c, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \coarse_time_0_r\);
    
    \counter_delta_snapshot_RNO_4[4]\ : NOR2A
      port map(A => N_384, B => \counter_delta_snapshot[4]_net_1\, 
        Y => counter_delta_snapshot_e4_i_a2_0);
    
    \counter_delta_snapshot_RNO_3[6]\ : NOR2A
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => counter_delta_snapshot_e6_i_a2_0, Y => N_455);
    
    counter_delta_snapshot_e27_0_0_o2_m6_e_1 : NOR2
      port map(A => \counter_delta_snapshot[19]_net_1\, B => 
        \counter_delta_snapshot[18]_net_1\, Y => 
        start_snapshot_f22_0_a2_11_0_a2_2_i);
    
    \counter_delta_f0[10]\ : DFN1E0C0
      port map(D => N_19, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9_0, Q => \counter_delta_f0[10]_net_1\);
    
    \counter_delta_snapshot_RNO_0[11]\ : OR3
      port map(A => N_391, B => \counter_delta_snapshot_i[11]\, C
         => N_504_0, Y => N_503);
    
    \counter_delta_f0_RNO[6]\ : MX2
      port map(A => delta_f2_f0(6), B => N_87_i_i, S => N_57, Y
         => N_11);
    
    start_snapshot_f22_0_a2 : NOR2
      port map(A => un12_start_snapshot_fothers_temp_NE, B => 
        start_snapshot_f22_0_a2_1, Y => N_7);
    
    \counter_delta_snapshot[5]\ : DFN1P0
      port map(D => N_376_i_0, CLK => HCLK_c, PRE => HRESETn_c, Q
         => \counter_delta_snapshot_i[5]\);
    
    \counter_delta_f0_RNO_0[12]\ : OAI1
      port map(A => N_67, B => \counter_delta_f0[11]_net_1\, C
         => counter_delta_f0_n12_0_0_a2_0, Y => N_252);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_14\ : XNOR2
      port map(A => \counter_delta_snapshot[13]_net_1\, B => 
        delta_snapshot(13), Y => N_133_i_i);
    
    \counter_delta_snapshot_RNO_3[4]\ : OR2B
      port map(A => counter_delta_snapshot_e4_i_a2_0, B => 
        \counter_delta_snapshot_RNIRV6E4[23]_net_1\, Y => N_445);
    
    \counter_delta_snapshot_RNO_2[18]\ : OR3
      port map(A => N_398, B => 
        \counter_delta_snapshot[18]_net_1\, C => N_504, Y => 
        N_176);
    
    \counter_delta_snapshot[0]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[0]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[0]_net_1\);
    
    \counter_delta_snapshot[7]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[7]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[7]_net_1\);
    
    \counter_delta_snapshot_RNO_1[13]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[13]_net_1\, C => N_285, Y => 
        counter_delta_snapshot_e13_i_0_0);
    
    start_snapshot_f1_RNO_1 : NOR3C
      port map(A => N_113_i_i_0, B => N_112_i_i_0, C => 
        start_snapshot_f12_0_a2_3, Y => start_snapshot_f12_0_a2_6);
    
    \counter_delta_f0_RNIGAGV2[24]\ : OR3
      port map(A => N_62, B => \counter_delta_f0[23]_net_1\, C
         => \counter_delta_f0[24]_net_1\, Y => N_66);
    
    \counter_delta_snapshot_RNO_2[9]\ : NOR3B
      port map(A => N_389, B => \counter_delta_snapshot[9]_net_1\, 
        C => N_504_0, Y => N_472);
    
    \counter_delta_f0_RNIPCA8[4]\ : NOR2
      port map(A => \counter_delta_f0[5]_net_1\, B => 
        \counter_delta_f0[4]_net_1\, Y => N_273);
    
    \counter_delta_f0_RNO[12]\ : AO1C
      port map(A => N_99, B => N_57_0, C => N_252, Y => 
        counter_delta_f0_n12);
    
    \counter_delta_snapshot[9]\ : DFN1C0
      port map(D => \counter_delta_snapshot_RNO[9]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_delta_snapshot[9]_net_1\);
    
    \counter_delta_snapshot_RNO_1[15]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[15]_net_1\, C => N_478, Y => 
        counter_delta_snapshot_e15_i_0_0);
    
    \counter_delta_snapshot_RNO[10]\ : NOR3
      port map(A => N_476, B => counter_delta_snapshot_e10_i_0, C
         => N_477, Y => \counter_delta_snapshot_RNO[10]_net_1\);
    
    \counter_delta_f0[11]\ : DFN1E0C0
      port map(D => N_275, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9_0, Q => \counter_delta_f0[11]_net_1\);
    
    \counter_delta_snapshot_RNO_0[22]\ : OR3C
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => \counter_delta_snapshot[22]_net_1\, C => N_402, Y
         => N_186);
    
    start_snapshot_f1_RNO_4 : XA1A
      port map(A => delta_f2_f1(9), B => 
        \counter_delta_f0[9]_net_1\, C => N_108_i_i_0, Y => 
        start_snapshot_f12_0_a2_4);
    
    \counter_delta_snapshot_RNO_0[12]\ : NOR2
      port map(A => N_505, B => delta_snapshot(12), Y => N_496);
    
    \counter_delta_snapshot_RNO[15]\ : NOR3
      port map(A => N_480, B => counter_delta_snapshot_e15_i_0_0, 
        C => N_482, Y => N_8);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_18\ : XNOR2
      port map(A => \counter_delta_snapshot[15]_net_1\, B => 
        delta_snapshot(15), Y => N_135_i_i);
    
    \counter_delta_snapshot_RNO_1[14]\ : AO1D
      port map(A => un2_coarse_time_0_0, B => 
        \counter_delta_snapshot[14]_net_1\, C => N_484, Y => 
        counter_delta_snapshot_e14_i_0_0);
    
    \counter_delta_f0_RNO_1[14]\ : NOR2B
      port map(A => \counter_delta_f0[14]_net_1\, B => N_57_0, Y
         => counter_delta_f0_n14_0_0_a2_0);
    
    \counter_delta_snapshot_RNO_0[19]\ : AOI1B
      port map(A => counter_delta_snapshot_e19_i_i_a2_0, B => 
        counter_delta_snapshot_e27_0_0_o2_N_7_0, C => N_178, Y
         => counter_delta_snapshot_e19_i_i_0);
    
    \counter_delta_f0[26]\ : DFN1E0C0
      port map(D => N_34, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_9, Q => \counter_delta_f0[26]_net_1\);
    
    \counter_delta_snapshot_RNO_4[6]\ : OR2A
      port map(A => N_386, B => \counter_delta_snapshot[6]_net_1\, 
        Y => counter_delta_snapshot_e6_i_a2_0);
    
    \counter_delta_snapshot_RNO[13]\ : NOR3
      port map(A => N_287, B => counter_delta_snapshot_e13_i_0_0, 
        C => N_288, Y => N_26);
    
    \counter_delta_snapshot_RNO_0[7]\ : NOR2
      port map(A => N_505, B => delta_snapshot(7), Y => N_462);
    
    \counter_delta_snapshot_RNO_0[26]\ : AO1B
      port map(A => \counter_delta_snapshot_RNIRV6E4[23]_net_1\, 
        B => N_406, C => un2_coarse_time_0, Y => 
        counter_delta_snapshot_e26_0_0_0_tz);
    
    \op_eq.un12_start_snapshot_fothers_temp_NE_RNO_16\ : XA1A
      port map(A => delta_snapshot(14), B => 
        \counter_delta_snapshot[14]_net_1\, C => N_135_i_i, Y => 
        un12_start_snapshot_fothers_temp_NE_3);
    
    \counter_delta_snapshot_RNO_0[16]\ : OA1A
      port map(A => \counter_delta_snapshot[16]_net_1\, B => 
        un2_coarse_time_0_0, C => N_168, Y => 
        counter_delta_snapshot_e16_i_i_0);
    
    start_snapshot_f1_RNO_3 : XA1A
      port map(A => delta_f2_f1(6), B => 
        \counter_delta_f0[6]_net_1\, C => N_82_i_i_0, Y => 
        start_snapshot_f12_0_a2_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\ is

    port( status_new_err    : out   std_logic_vector(3 to 3);
          valid_ack         : in    std_logic_vector(3 to 3);
          valid_out         : out   std_logic_vector(3 to 3);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f3_out_valid : in    std_logic
        );

end 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\ is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal state_1_sqmuxa_1_i, N_6_i_i_0, \valid_out[3]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    valid_out(3) <= \valid_out[3]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    error : DFN1C0
      port map(D => state_1_sqmuxa_1_i, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => status_new_err(3));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state[0]\ : DFN1C0
      port map(D => N_6_i_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => \valid_out[3]\);
    
    error_RNO : NOR3B
      port map(A => \valid_out[3]\, B => data_f3_out_valid, C => 
        valid_ack(3), Y => state_1_sqmuxa_1_i);
    
    \state_RNO[0]\ : AX1
      port map(A => valid_ack(3), B => \valid_out[3]\, C => 
        data_f3_out_valid, Y => N_6_i_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\ is

    port( status_new_err    : out   std_logic_vector(1 to 1);
          valid_out_i       : out   std_logic_vector(1 to 1);
          valid_ack         : in    std_logic_vector(1 to 1);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f1_out_valid : in    std_logic
        );

end 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\ is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal state_1_sqmuxa_1, N_6_i_i_0, \valid_out_i[1]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    valid_out_i(1) <= \valid_out_i[1]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    error : DFN1C0
      port map(D => state_1_sqmuxa_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => status_new_err(1));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state[0]\ : DFN1P0
      port map(D => N_6_i_i_0, CLK => HCLK_c, PRE => HRESETn_c, Q
         => \valid_out_i[1]\);
    
    error_RNO : NOR3A
      port map(A => data_f1_out_valid, B => valid_ack(1), C => 
        \valid_out_i[1]\, Y => state_1_sqmuxa_1);
    
    \state_RNO[0]\ : AX1D
      port map(A => valid_ack(1), B => \valid_out_i[1]\, C => 
        data_f1_out_valid, Y => N_6_i_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_burst is

    port( sample_f3_wdata   : in    std_logic_vector(95 downto 0);
          data_f3_out       : out   std_logic_vector(159 downto 64);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f3_out_valid : out   std_logic;
          enable_f3         : in    std_logic;
          sample_f3_val     : in    std_logic
        );

end lpp_waveform_burst;

architecture DEF_ARCH of lpp_waveform_burst is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal data_out_valid_3, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \data_out[91]\ : DFN1C0
      port map(D => sample_f3_wdata(27), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(91));
    
    \data_out[124]\ : DFN1C0
      port map(D => sample_f3_wdata(60), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(124));
    
    \data_out[120]\ : DFN1C0
      port map(D => sample_f3_wdata(56), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(120));
    
    \data_out[138]\ : DFN1C0
      port map(D => sample_f3_wdata(74), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(138));
    
    \data_out[105]\ : DFN1C0
      port map(D => sample_f3_wdata(41), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(105));
    
    \data_out[126]\ : DFN1C0
      port map(D => sample_f3_wdata(62), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(126));
    
    \data_out[74]\ : DFN1C0
      port map(D => sample_f3_wdata(10), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(74));
    
    \data_out[154]\ : DFN1C0
      port map(D => sample_f3_wdata(90), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(154));
    
    \data_out[150]\ : DFN1C0
      port map(D => sample_f3_wdata(86), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(150));
    
    \data_out[102]\ : DFN1C0
      port map(D => sample_f3_wdata(38), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(102));
    
    \data_out[156]\ : DFN1C0
      port map(D => sample_f3_wdata(92), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(156));
    
    \data_out[93]\ : DFN1C0
      port map(D => sample_f3_wdata(29), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(93));
    
    \data_out[128]\ : DFN1C0
      port map(D => sample_f3_wdata(64), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(128));
    
    data_out_valid : DFN1C0
      port map(D => data_out_valid_3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out_valid);
    
    \data_out[69]\ : DFN1C0
      port map(D => sample_f3_wdata(5), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(69));
    
    \data_out[141]\ : DFN1C0
      port map(D => sample_f3_wdata(77), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(141));
    
    \data_out[99]\ : DFN1C0
      port map(D => sample_f3_wdata(35), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(99));
    
    \data_out[147]\ : DFN1C0
      port map(D => sample_f3_wdata(83), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(147));
    
    \data_out[87]\ : DFN1C0
      port map(D => sample_f3_wdata(23), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(87));
    
    \data_out[149]\ : DFN1C0
      port map(D => sample_f3_wdata(85), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(149));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \data_out[86]\ : DFN1C0
      port map(D => sample_f3_wdata(22), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(86));
    
    \data_out[158]\ : DFN1C0
      port map(D => sample_f3_wdata(94), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(158));
    
    \data_out[113]\ : DFN1C0
      port map(D => sample_f3_wdata(49), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(113));
    
    \data_out[65]\ : DFN1C0
      port map(D => sample_f3_wdata(1), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(65));
    
    \data_out[95]\ : DFN1C0
      port map(D => sample_f3_wdata(31), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(95));
    
    \data_out[92]\ : DFN1C0
      port map(D => sample_f3_wdata(28), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(92));
    
    \data_out[77]\ : DFN1C0
      port map(D => sample_f3_wdata(13), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(77));
    
    \data_out[145]\ : DFN1C0
      port map(D => sample_f3_wdata(81), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(145));
    
    \data_out[131]\ : DFN1C0
      port map(D => sample_f3_wdata(67), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(131));
    
    \data_out[76]\ : DFN1C0
      port map(D => sample_f3_wdata(12), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(76));
    
    \data_out[137]\ : DFN1C0
      port map(D => sample_f3_wdata(73), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(137));
    
    \data_out[139]\ : DFN1C0
      port map(D => sample_f3_wdata(75), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(139));
    
    \data_out[114]\ : DFN1C0
      port map(D => sample_f3_wdata(50), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(114));
    
    \data_out[80]\ : DFN1C0
      port map(D => sample_f3_wdata(16), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(80));
    
    \data_out[64]\ : DFN1C0
      port map(D => sample_f3_wdata(0), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(64));
    
    \data_out[110]\ : DFN1C0
      port map(D => sample_f3_wdata(46), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(110));
    
    \data_out[103]\ : DFN1C0
      port map(D => sample_f3_wdata(39), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(103));
    
    \data_out[142]\ : DFN1C0
      port map(D => sample_f3_wdata(78), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(142));
    
    \data_out[94]\ : DFN1C0
      port map(D => sample_f3_wdata(30), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(94));
    
    \data_out[88]\ : DFN1C0
      port map(D => sample_f3_wdata(24), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(88));
    
    \data_out[116]\ : DFN1C0
      port map(D => sample_f3_wdata(52), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(116));
    
    \data_out[121]\ : DFN1C0
      port map(D => sample_f3_wdata(57), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(121));
    
    \data_out[127]\ : DFN1C0
      port map(D => sample_f3_wdata(63), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(127));
    
    \data_out[129]\ : DFN1C0
      port map(D => sample_f3_wdata(65), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(129));
    
    \data_out[135]\ : DFN1C0
      port map(D => sample_f3_wdata(71), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(135));
    
    \data_out[70]\ : DFN1C0
      port map(D => sample_f3_wdata(6), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(70));
    
    data_out_valid_RNO : NOR2B
      port map(A => sample_f3_val, B => enable_f3, Y => 
        data_out_valid_3);
    
    \data_out[118]\ : DFN1C0
      port map(D => sample_f3_wdata(54), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(118));
    
    \data_out[104]\ : DFN1C0
      port map(D => sample_f3_wdata(40), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(104));
    
    \data_out[100]\ : DFN1C0
      port map(D => sample_f3_wdata(36), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(100));
    
    \data_out[78]\ : DFN1C0
      port map(D => sample_f3_wdata(14), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(78));
    
    \data_out[151]\ : DFN1C0
      port map(D => sample_f3_wdata(87), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(151));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \data_out[157]\ : DFN1C0
      port map(D => sample_f3_wdata(93), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(157));
    
    \data_out[106]\ : DFN1C0
      port map(D => sample_f3_wdata(42), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(106));
    
    \data_out[159]\ : DFN1C0
      port map(D => sample_f3_wdata(95), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(159));
    
    \data_out[132]\ : DFN1C0
      port map(D => sample_f3_wdata(68), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(132));
    
    \data_out[125]\ : DFN1C0
      port map(D => sample_f3_wdata(61), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(125));
    
    \data_out[67]\ : DFN1C0
      port map(D => sample_f3_wdata(3), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(67));
    
    \data_out[81]\ : DFN1C0
      port map(D => sample_f3_wdata(17), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(81));
    
    \data_out[97]\ : DFN1C0
      port map(D => sample_f3_wdata(33), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(97));
    
    \data_out[66]\ : DFN1C0
      port map(D => sample_f3_wdata(2), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(66));
    
    \data_out[108]\ : DFN1C0
      port map(D => sample_f3_wdata(44), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(108));
    
    \data_out[96]\ : DFN1C0
      port map(D => sample_f3_wdata(32), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(96));
    
    \data_out[143]\ : DFN1C0
      port map(D => sample_f3_wdata(79), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(143));
    
    \data_out[122]\ : DFN1C0
      port map(D => sample_f3_wdata(58), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(122));
    
    \data_out[155]\ : DFN1C0
      port map(D => sample_f3_wdata(91), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(155));
    
    \data_out[71]\ : DFN1C0
      port map(D => sample_f3_wdata(7), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(71));
    
    \data_out[152]\ : DFN1C0
      port map(D => sample_f3_wdata(88), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(152));
    
    \data_out[83]\ : DFN1C0
      port map(D => sample_f3_wdata(19), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(83));
    
    \data_out[144]\ : DFN1C0
      port map(D => sample_f3_wdata(80), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(144));
    
    \data_out[140]\ : DFN1C0
      port map(D => sample_f3_wdata(76), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(140));
    
    \data_out[111]\ : DFN1C0
      port map(D => sample_f3_wdata(47), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(111));
    
    \data_out[90]\ : DFN1C0
      port map(D => sample_f3_wdata(26), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(90));
    
    \data_out[89]\ : DFN1C0
      port map(D => sample_f3_wdata(25), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(89));
    
    \data_out[68]\ : DFN1C0
      port map(D => sample_f3_wdata(4), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(68));
    
    \data_out[117]\ : DFN1C0
      port map(D => sample_f3_wdata(53), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(117));
    
    \data_out[146]\ : DFN1C0
      port map(D => sample_f3_wdata(82), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(146));
    
    \data_out[133]\ : DFN1C0
      port map(D => sample_f3_wdata(69), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(133));
    
    \data_out[119]\ : DFN1C0
      port map(D => sample_f3_wdata(55), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(119));
    
    \data_out[98]\ : DFN1C0
      port map(D => sample_f3_wdata(34), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(98));
    
    \data_out[73]\ : DFN1C0
      port map(D => sample_f3_wdata(9), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(73));
    
    \data_out[85]\ : DFN1C0
      port map(D => sample_f3_wdata(21), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(85));
    
    \data_out[82]\ : DFN1C0
      port map(D => sample_f3_wdata(18), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(82));
    
    \data_out[79]\ : DFN1C0
      port map(D => sample_f3_wdata(15), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(79));
    
    \data_out[148]\ : DFN1C0
      port map(D => sample_f3_wdata(84), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(148));
    
    \data_out[123]\ : DFN1C0
      port map(D => sample_f3_wdata(59), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(123));
    
    \data_out[101]\ : DFN1C0
      port map(D => sample_f3_wdata(37), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(101));
    
    \data_out[134]\ : DFN1C0
      port map(D => sample_f3_wdata(70), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(134));
    
    \data_out[115]\ : DFN1C0
      port map(D => sample_f3_wdata(51), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(115));
    
    \data_out[130]\ : DFN1C0
      port map(D => sample_f3_wdata(66), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(130));
    
    \data_out[107]\ : DFN1C0
      port map(D => sample_f3_wdata(43), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(107));
    
    \data_out[109]\ : DFN1C0
      port map(D => sample_f3_wdata(45), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(109));
    
    \data_out[136]\ : DFN1C0
      port map(D => sample_f3_wdata(72), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(136));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \data_out[84]\ : DFN1C0
      port map(D => sample_f3_wdata(20), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(84));
    
    \data_out[75]\ : DFN1C0
      port map(D => sample_f3_wdata(11), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(75));
    
    \data_out[72]\ : DFN1C0
      port map(D => sample_f3_wdata(8), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(72));
    
    \data_out[153]\ : DFN1C0
      port map(D => sample_f3_wdata(89), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(153));
    
    \data_out[112]\ : DFN1C0
      port map(D => sample_f3_wdata(48), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f3_out(112));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\ is

    port( status_new_err    : out   std_logic_vector(2 to 2);
          valid_ack         : in    std_logic_vector(2 to 2);
          valid_out         : out   std_logic_vector(2 to 2);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f2_out_valid : in    std_logic
        );

end 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\ is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal state_1_sqmuxa_1, N_6_i_i_0, \valid_out[2]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    valid_out(2) <= \valid_out[2]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    error : DFN1C0
      port map(D => state_1_sqmuxa_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => status_new_err(2));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state[0]\ : DFN1C0
      port map(D => N_6_i_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => \valid_out[2]\);
    
    error_RNO : NOR3B
      port map(A => \valid_out[2]\, B => data_f2_out_valid, C => 
        valid_ack(2), Y => state_1_sqmuxa_1);
    
    \state_RNO[0]\ : AX1
      port map(A => valid_ack(2), B => \valid_out[2]\, C => 
        data_f2_out_valid, Y => N_6_i_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\ is

    port( status_new_err    : out   std_logic_vector(0 to 0);
          valid_ack         : in    std_logic_vector(0 to 0);
          valid_out         : out   std_logic_vector(0 to 0);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f0_out_valid : in    std_logic
        );

end 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\ is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal state_1_sqmuxa_1, N_6_i_i_0, \valid_out[0]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    valid_out(0) <= \valid_out[0]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    error : DFN1C0
      port map(D => state_1_sqmuxa_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => status_new_err(0));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state[0]\ : DFN1C0
      port map(D => N_6_i_i_0, CLK => HCLK_c, CLR => HRESETn_c, Q
         => \valid_out[0]\);
    
    error_RNO : NOR3B
      port map(A => \valid_out[0]\, B => data_f0_out_valid, C => 
        valid_ack(0), Y => state_1_sqmuxa_1);
    
    \state_RNO[0]\ : AX1
      port map(A => valid_ack(0), B => \valid_out[0]\, C => 
        data_f0_out_valid, Y => N_6_i_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ1 is

    port( ready_i_0             : out   std_logic_vector(1 to 1);
          Raddr_vect_RNICA1PH   : out   std_logic_vector(1 to 1);
          data_mem_wen_i_0      : inout std_logic_vector(2 downto 1) := (others => 'Z');
          Raddr_vect_RNIIMQ5I   : out   std_logic_vector(4 to 4);
          Raddr_vect_RNIE6Q5I   : out   std_logic_vector(3 to 3);
          Raddr_vect_RNIKA2PH   : out   std_logic_vector(2 to 2);
          data_addr_r_iv_i_3    : in    std_logic_vector(4 downto 0);
          Raddr_vect_RNI4A0PH   : out   std_logic_vector(0 to 0);
          data_addr_r_iv_i_a2_2 : in    std_logic_vector(4 to 4);
          data_wen              : in    std_logic_vector(1 to 1);
          data_mem_ren_i_0      : inout std_logic_vector(1 downto 0) := (others => 'Z');
          data_ren              : in    std_logic_vector(1 to 1);
          data_ren_1z           : in    std_logic;
          HRESETn_c             : in    std_logic;
          HCLK_c                : in    std_logic;
          N_166                 : out   std_logic;
          N_126                 : out   std_logic;
          N_150                 : out   std_logic;
          N_134                 : out   std_logic;
          N_142                 : out   std_logic;
          N_165                 : in    std_logic;
          N_158                 : out   std_logic;
          un20_time_write       : in    std_logic;
          N_68                  : in    std_logic;
          N_164                 : in    std_logic;
          N_120_i               : out   std_logic;
          N_44                  : in    std_logic;
          N_52                  : in    std_logic;
          N_60                  : in    std_logic;
          N_76                  : in    std_logic;
          N_86                  : out   std_logic;
          N_75                  : in    std_logic;
          N_59                  : in    std_logic;
          N_51                  : in    std_logic;
          N_43                  : in    std_logic;
          N_67                  : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ1;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ1 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_12, \data_mem_addr_w_1[1]\, \data_mem_addr_w_1[0]\, 
        N_4, \data_mem_addr_w_1[3]\, \DWACT_FINC_E[0]\, N_12_0, 
        \data_mem_addr_r_1[1]\, \data_mem_addr_r_1[0]\, N_4_0, 
        \data_mem_addr_r_1[3]\, \DWACT_FINC_E_0[0]\, 
        \un26_sfull_s\, \un26_sfull_s_tz\, \sFull\, un5_sfull_s_4, 
        \data_addr_r_iv_i_4[1]\, \data_addr_r_iv_i_4[4]\, 
        \data_mem_addr_r_1[4]\, \data_addr_r_iv_i_4[3]\, 
        \data_addr_r_iv_i_4[2]\, \data_mem_addr_r_1[2]\, 
        \data_addr_r_iv_i_4[0]\, \data_addr_r_iv_i_a2_3[4]\, 
        un7_sempty_s_4, un7_sempty_s_1, un7_sempty_s_0, 
        un7_sempty_s_2, \un10_raddr_vect_s[3]\, sEmpty_RNO_7_0, 
        \un10_raddr_vect_s[1]\, sEmpty_RNO_6_2, 
        \un10_raddr_vect_s[0]\, un5_sfull_s_4_2, 
        \un8_waddr_vect_s[3]\, \un26_sfull_s_tz_RNO_7\, 
        un5_sfull_s_4_1, \un8_waddr_vect_s[1]\, 
        \un26_sfull_s_tz_RNO_4\, un5_sfull_s_4_0, 
        \un8_waddr_vect_s[0]\, ADD_5x5_fast_I11_Y_i_a2_0, 
        \data_mem_addr_w_1[2]\, N_109, ADD_5x5_fast_I11_Y_0, 
        N_89_i, N80, SUM2_0_0, ADD_5x5_fast_I11_un1_Y_0, N81, 
        N_85_i, N_105_1, ADD_7x7_fast_I19_Y_i_o4_1_0, N_87, 
        un1_waddr_vect_slto3_0, un2_raddr_vect_slto3_0, 
        un1_waddr_vect_slt4, \un60_ready1[4]\, CO1_tz, N_12_1, 
        N_17, N_18, I11_un1_Y, un7_sempty_s, Waddr_vect_n4, 
        \data_mem_addr_w_1[4]\, Waddr_vect_14_0, Waddr_vect_c2, 
        Waddr_vect_n2, un1_waddr_vect_s, Waddr_vect_n2_tz, 
        Waddr_vect_n3, N_9, N165, N_14_1, N_23, N_75_i_0, 
        \un75_ready1[4]\, ADD_5x5_fast_I8_un1_Y_0, 
        \un75_ready0_1[4]\, \un60_ready0[4]\, N_13, 
        \un75_ready0[4]\, un62_readylto4, un77_ready, un69_ready, 
        N_198, N107, N161, N_197, \un75_ready1[5]\, N_16_i_i_0, 
        N_196, N83, un2_raddr_vect_slto1, un2_raddr_vect_s, 
        Waddr_vect_e0, Waddr_vect_e1, Waddr_vect_n1_i, 
        Waddr_vect_e4, Waddr_vect_e2, I_20_9, I_9_17, 
        \un10_raddr_vect_s[4]\, \un10_raddr_vect_s[2]\, 
        Waddr_vect_e3, I_13_17, I_5_17, I_20_10, I_13_18, I_9_18, 
        I_5_18, sEmpty_RNO_11, un1_sempty_s, \sEmpty\, N_9_0, 
        N_13_0, N_12_2, N_11, N_8, N_10, N_9_1, N_7, N_4_1, N_5, 
        N_6, N_9_2, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    sFull : DFN1C0
      port map(D => \un26_sfull_s\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \Raddr_vect_RNICA1PH[1]\ : NOR3C
      port map(A => \data_addr_r_iv_i_4[1]\, B => 
        data_addr_r_iv_i_3(1), C => N_68, Y => 
        Raddr_vect_RNICA1PH(1));
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => data_mem_wen_i_0(1), C
         => \data_mem_addr_w_1[0]\, Y => Waddr_vect_e0);
    
    \Raddr_vect_RNIA2FB1[0]\ : MX2
      port map(A => \un60_ready1[4]\, B => \un60_ready0[4]\, S
         => \data_mem_addr_r_1[0]\, Y => un62_readylto4);
    
    un75_ready_1_16_ADD_5x5_fast_I8_un1_Y : NOR3A
      port map(A => N81, B => N_85_i, C => N_105_1, Y => 
        ADD_5x5_fast_I8_un1_Y_0);
    
    \Raddr_vect_RNI7873[3]\ : XNOR2
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \data_mem_addr_r_1[3]\, Y => N_87);
    
    \Waddr_vect_RNIIOD6[0]\ : AO1B
      port map(A => \data_mem_addr_w_1[1]\, B => 
        \data_mem_addr_w_1[0]\, C => un1_waddr_vect_slto3_0, Y
         => un1_waddr_vect_slt4);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_1[0]\);
    
    sEmpty_RNIANF32 : NOR3A
      port map(A => data_ren_1z, B => un20_time_write, C => 
        \sEmpty\, Y => data_mem_ren_i_0(1));
    
    \Waddr_vect_RNO[3]\ : MX2A
      port map(A => Waddr_vect_n3, B => \data_mem_addr_w_1[3]\, S
         => data_mem_wen_i_0(1), Y => Waddr_vect_e3);
    
    un26_sfull_s_tz_RNO_5 : OR2A
      port map(A => un1_waddr_vect_s, B => \data_mem_addr_w_1[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    \Raddr_vect_RNI3O63[1]\ : NOR2A
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \data_mem_addr_w_1[1]\, Y => N_105_1);
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \data_mem_addr_r_1[0]\, Y => N_12_0);
    
    un26_sfull_s_tz_RNO_3 : OR2B
      port map(A => I_5_17, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[1]\);
    
    \ready_gen.un69_ready_0_I_8\ : OR2A
      port map(A => \data_mem_addr_w_1[4]\, B => 
        \data_mem_addr_r_1[4]\, Y => N_11);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \data_mem_addr_w_1[1]\, Y => I_5_17);
    
    sEmpty_RNO_0 : NOR3B
      port map(A => data_ren_1z, B => un7_sempty_s_4, C => 
        un20_time_write, Y => un7_sempty_s);
    
    \Waddr_vect_RNIE4CV[3]\ : OR3A
      port map(A => N_165, B => data_mem_wen_i_0(1), C => 
        \data_mem_addr_w_1[3]\, Y => N_134);
    
    un60_ready_1_1_0_SUM2_0 : AX1C
      port map(A => N_87, B => CO1_tz, C => SUM2_0_0, Y => 
        \un60_ready1[4]\);
    
    \Raddr_vect_RNIU7FE[4]\ : NOR2B
      port map(A => I_13_18, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    un26_sfull_s_tz_RNO_6 : OR2B
      port map(A => I_13_17, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    \Raddr_vect_RNI0G18[4]\ : AO1B
      port map(A => un2_raddr_vect_slto3_0, B => 
        un2_raddr_vect_slto1, C => \data_mem_addr_r_1[4]\, Y => 
        un2_raddr_vect_s);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_r_1[0]\, B => 
        \data_mem_addr_r_1[1]\, C => \data_mem_addr_r_1[2]\, Y
         => N_9_0);
    
    \Raddr_vect_RNIB44A2[0]\ : MX2C
      port map(A => N107, B => N161, S => \data_mem_addr_r_1[0]\, 
        Y => N_198);
    
    \ready_gen.un69_ready_0_I_2\ : OR2A
      port map(A => \data_mem_addr_w_1[2]\, B => 
        \data_mem_addr_r_1[2]\, Y => N_5);
    
    \ready_gen.un69_ready_0_I_7\ : AO1C
      port map(A => \data_mem_addr_w_1[2]\, B => 
        \data_mem_addr_r_1[2]\, C => N_4_1, Y => N_10);
    
    \Raddr_vect_RNIK66A4[1]\ : OA1A
      port map(A => data_mem_ren_i_0(1), B => 
        \data_mem_addr_r_1[1]\, C => N_67, Y => 
        \data_addr_r_iv_i_4[1]\);
    
    \Waddr_vect_RNO[4]\ : MX2A
      port map(A => Waddr_vect_n4, B => \data_mem_addr_w_1[4]\, S
         => data_mem_wen_i_0(1), Y => Waddr_vect_e4);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_1[1]\);
    
    un75_ready_0_0_0_ADD_7x7_fast_I32_Y_0 : XOR2
      port map(A => N165, B => \un75_ready0_1[4]\, Y => 
        \un75_ready0[4]\);
    
    un60_ready_0_0_0_ADD_5x5_fast_I9_Y_i_o2 : AO13
      port map(A => \data_mem_addr_w_1[1]\, B => 
        \data_mem_addr_w_1[0]\, C => \data_mem_addr_r_1[1]\, Y
         => N_9);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_9_2, B => \data_mem_addr_w_1[3]\, Y => 
        I_13_17);
    
    sFull_RNI8GOT : OR2B
      port map(A => data_mem_wen_i_0(1), B => N_165, Y => N_166);
    
    GND_i : GND
      port map(Y => \GND\);
    
    sEmpty_RNO_7 : XNOR2
      port map(A => \un10_raddr_vect_s[4]\, B => 
        \data_mem_addr_w_1[4]\, Y => sEmpty_RNO_7_0);
    
    sEmpty_RNIGNUI8 : NOR2B
      port map(A => \data_addr_r_iv_i_a2_3[4]\, B => 
        data_addr_r_iv_i_a2_2(4), Y => N_86);
    
    \Raddr_vect_RNIT38B[4]\ : NOR2B
      port map(A => I_5_18, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[1]\);
    
    un26_sfull_s_tz_RNO_0 : XA1
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \un8_waddr_vect_s[1]\, C => \un26_sfull_s_tz_RNO_4\, Y
         => un5_sfull_s_4_1);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \data_mem_addr_w_1[1]\, C => \data_mem_addr_w_1[2]\, Y
         => N_9_2);
    
    \Raddr_vect_RNI5073[2]\ : XNOR2
      port map(A => \data_mem_addr_w_1[2]\, B => 
        \data_mem_addr_r_1[2]\, Y => N_85_i);
    
    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \data_mem_addr_w_1[1]\, B => 
        \data_mem_addr_w_1[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    \Raddr_vect[2]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => data_mem_ren_i_0(1), Q => 
        \data_mem_addr_r_1[2]\);
    
    un60_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0 : OR2A
      port map(A => \data_mem_addr_r_1[3]\, B => 
        \data_mem_addr_w_1[3]\, Y => N_13);
    
    sEmpty_RNIJEV64 : NOR2
      port map(A => data_mem_ren_i_0(1), B => data_mem_ren_i_0(0), 
        Y => \data_addr_r_iv_i_a2_3[4]\);
    
    \ready_gen.un69_ready_0_I_4\ : OR2A
      port map(A => \data_mem_addr_r_1[4]\, B => 
        \data_mem_addr_w_1[4]\, Y => N_7);
    
    un75_ready_1_16_ADD_5x5_fast_I1_P0N : OR2A
      port map(A => \data_mem_addr_r_1[2]\, B => N_87, Y => N81);
    
    un75_ready_0_0_0_ADD_7x7_fast_I23_Y_0_o2_1 : OA1C
      port map(A => N165, B => N_89_i, C => N_23, Y => N_14_1);
    
    un60_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3_0 : NOR2B
      port map(A => N_9, B => \data_mem_addr_w_1[2]\, Y => N_18);
    
    \Waddr_vect_RNO_0[4]\ : AXO1
      port map(A => un1_waddr_vect_slt4, B => 
        \data_mem_addr_w_1[4]\, C => Waddr_vect_14_0, Y => 
        Waddr_vect_n4);
    
    sFull_RNIBVR9 : OR2
      port map(A => \sFull\, B => data_wen(1), Y => 
        data_mem_wen_i_0(1));
    
    \Raddr_vect_RNIT3LC6[0]\ : AOI1
      port map(A => N_197, B => N_196, C => N_198, Y => 
        un77_ready);
    
    \Raddr_vect_RNI9G73_0[4]\ : NOR2A
      port map(A => \data_mem_addr_r_1[4]\, B => 
        \data_mem_addr_w_1[4]\, Y => N_75_i_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un75_ready_0_0_0_ADD_7x7_fast_I23_Y_0 : OR2B
      port map(A => N_14_1, B => N_75_i_0, Y => N161);
    
    un75_ready_1_16_ADD_5x5_fast_I2_G0N : OR2
      port map(A => N_109, B => N_89_i, Y => N83);
    
    sEmpty_RNO : OR2
      port map(A => un7_sempty_s, B => un1_sempty_s, Y => 
        sEmpty_RNO_11);
    
    \Waddr_vect[3]\ : DFN1C0
      port map(D => Waddr_vect_e3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_1[3]\);
    
    un26_sfull_s : AND2
      port map(A => data_ren(1), B => \un26_sfull_s_tz\, Y => 
        \un26_sfull_s\);
    
    \Waddr_vect_RNIB473[3]\ : NOR2
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \data_mem_addr_w_1[2]\, Y => un1_waddr_vect_slto3_0);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_w_1[1]\, B => 
        \data_mem_addr_w_1[0]\, Y => N_12);
    
    sEmpty_RNO_3 : XA1A
      port map(A => \data_mem_addr_w_1[1]\, B => 
        \un10_raddr_vect_s[1]\, C => sEmpty_RNO_6_2, Y => 
        un7_sempty_s_1);
    
    un26_sfull_s_tz_RNO_4 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_17, C => 
        \data_mem_addr_r_1[2]\, Y => \un26_sfull_s_tz_RNO_4\);
    
    un75_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4 : AO1B
      port map(A => ADD_7x7_fast_I19_Y_i_o4_1_0, B => N_9, C => 
        N80, Y => N165);
    
    un6_waddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \DWACT_FINC_E[0]\, Y => N_4);
    
    \Waddr_vect[4]\ : DFN1C0
      port map(D => Waddr_vect_e4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_1[4]\);
    
    \ready_gen.un69_ready_0_I_5\ : AO1C
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \data_mem_addr_w_1[1]\, C => N_6, Y => N_8);
    
    \Raddr_vect_RNIOM6A4[3]\ : OA1A
      port map(A => data_mem_ren_i_0(1), B => 
        \data_mem_addr_r_1[3]\, C => N_51, Y => 
        \data_addr_r_iv_i_4[3]\);
    
    \Raddr_vect_RNIE6Q5I[3]\ : NOR3C
      port map(A => \data_addr_r_iv_i_4[3]\, B => 
        data_addr_r_iv_i_3(3), C => N_52, Y => 
        Raddr_vect_RNIE6Q5I(3));
    
    \Waddr_vect_RNO_0[2]\ : OR2B
      port map(A => un1_waddr_vect_s, B => Waddr_vect_n2_tz, Y
         => Waddr_vect_n2);
    
    \Raddr_vect_RNI003G[4]\ : NOR2B
      port map(A => I_20_10, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[4]\);
    
    un75_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1_0 : AXOI5
      port map(A => N_87, B => \data_mem_addr_r_1[2]\, C => 
        \data_mem_addr_w_1[2]\, Y => ADD_7x7_fast_I19_Y_i_o4_1_0);
    
    \ready_gen.un69_ready_0_I_9\ : AO1C
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \data_mem_addr_r_1[3]\, C => N_7, Y => N_12_2);
    
    un26_sfull_s_tz : OR2
      port map(A => \sFull\, B => un5_sfull_s_4, Y => 
        \un26_sfull_s_tz\);
    
    un75_ready_0_0_0_ADD_7x7_fast_I33_Y_0_i_x2 : AX1E
      port map(A => N_14_1, B => N83, C => N_75_i_0, Y => 
        N_16_i_i_0);
    
    \Waddr_vect_RNID0CV[2]\ : OR3A
      port map(A => N_165, B => data_mem_wen_i_0(1), C => 
        \data_mem_addr_w_1[2]\, Y => N_142);
    
    \Raddr_vect_RNIKA2PH[2]\ : NOR3C
      port map(A => \data_addr_r_iv_i_4[2]\, B => 
        data_addr_r_iv_i_3(2), C => N_60, Y => 
        Raddr_vect_RNIKA2PH(2));
    
    \Raddr_vect_RNIUNK9[0]\ : NOR2A
      port map(A => un2_raddr_vect_s, B => \data_mem_addr_r_1[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    \Raddr_vect[0]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => data_mem_ren_i_0(1), Q => 
        \data_mem_addr_r_1[0]\);
    
    \Waddr_vect_RNO_0[3]\ : XAI1
      port map(A => \data_mem_addr_w_1[3]\, B => Waddr_vect_c2, C
         => un1_waddr_vect_s, Y => Waddr_vect_n3);
    
    \Raddr_vect_RNI9G73[4]\ : XNOR2
      port map(A => \data_mem_addr_w_1[4]\, B => 
        \data_mem_addr_r_1[4]\, Y => N_89_i);
    
    \Waddr_vect_RNIF8CV[4]\ : OR3A
      port map(A => N_165, B => data_mem_wen_i_0(1), C => 
        \data_mem_addr_w_1[4]\, Y => N_126);
    
    \Raddr_vect_RNIIU5A4[0]\ : OA1A
      port map(A => data_mem_ren_i_0(1), B => 
        \data_mem_addr_r_1[0]\, C => N_75, Y => 
        \data_addr_r_iv_i_4[0]\);
    
    \Raddr_vect_RNION3L8[0]\ : MX2
      port map(A => un62_readylto4, B => un77_ready, S => 
        un69_ready, Y => ready_i_0(1));
    
    un60_ready_1_1_0_SUM2_0_0 : XNOR2
      port map(A => N_109, B => N_89_i, Y => SUM2_0_0);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_12_0, B => \data_mem_addr_r_1[2]\, Y => 
        I_9_18);
    
    \ready_gen.un69_ready_0_I_1\ : OR2A
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \data_mem_addr_w_1[1]\, Y => N_4_1);
    
    \Raddr_vect_RNITJ63[1]\ : OR2B
      port map(A => \data_mem_addr_r_1[1]\, B => 
        \data_mem_addr_r_1[0]\, Y => un2_raddr_vect_slto1);
    
    un75_ready_0_0_0_ADD_7x7_fast_I32_Y_0_1 : XOR2
      port map(A => N_109, B => N_89_i, Y => \un75_ready0_1[4]\);
    
    un60_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2 : OR3
      port map(A => N_17, B => ADD_5x5_fast_I11_Y_i_a2_0, C => 
        N_18, Y => N_12_1);
    
    un75_ready_1_16_ADD_5x5_fast_I10_Y : OR3A
      port map(A => N_75_i_0, B => I11_un1_Y, C => 
        ADD_5x5_fast_I11_Y_0, Y => N107);
    
    \Waddr_vect_RNICSBV[1]\ : OR3A
      port map(A => N_165, B => data_mem_wen_i_0(1), C => 
        \data_mem_addr_w_1[1]\, Y => N_150);
    
    un75_ready_0_0_0_ADD_7x7_fast_I23_Y_0_a4 : NOR3B
      port map(A => N_9, B => ADD_7x7_fast_I19_Y_i_o4_1_0, C => 
        N_109, Y => N_23);
    
    un26_sfull_s_tz_RNO : NOR3C
      port map(A => un5_sfull_s_4_1, B => un5_sfull_s_4_0, C => 
        un5_sfull_s_4_2, Y => un5_sfull_s_4);
    
    un8_raddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_r_1[0]\, B => 
        \data_mem_addr_r_1[1]\, C => \data_mem_addr_r_1[2]\, Y
         => \DWACT_FINC_E_0[0]\);
    
    \Raddr_vect_RNIN2UH1[0]\ : MX2C
      port map(A => \un75_ready1[4]\, B => \un75_ready0[4]\, S
         => \data_mem_addr_r_1[0]\, Y => N_196);
    
    \Waddr_vect_RNIC4Q4[0]\ : NOR3C
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \data_mem_addr_w_1[1]\, C => \data_mem_addr_w_1[2]\, Y
         => Waddr_vect_c2);
    
    \Waddr_vect_RNO_1[4]\ : OR2B
      port map(A => Waddr_vect_c2, B => \data_mem_addr_w_1[3]\, Y
         => Waddr_vect_14_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Waddr_vect_RNIPG18[4]\ : OR2B
      port map(A => un1_waddr_vect_slt4, B => 
        \data_mem_addr_w_1[4]\, Y => un1_waddr_vect_s);
    
    un75_ready_1_16_ADD_5x5_fast_I11_un1_Y_0 : NOR3A
      port map(A => N81, B => N_85_i, C => N_105_1, Y => 
        ADD_5x5_fast_I11_un1_Y_0);
    
    un26_sfull_s_tz_RNO_7 : AX1E
      port map(A => un1_waddr_vect_s, B => I_20_9, C => 
        \data_mem_addr_r_1[4]\, Y => \un26_sfull_s_tz_RNO_7\);
    
    un6_waddr_vect_s_I_20 : XOR2
      port map(A => N_4, B => \data_mem_addr_w_1[4]\, Y => I_20_9);
    
    \Raddr_vect[1]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => data_mem_ren_i_0(1), Q => 
        \data_mem_addr_r_1[1]\);
    
    sEmpty_RNO_6 : XNOR2
      port map(A => \un10_raddr_vect_s[2]\, B => 
        \data_mem_addr_w_1[2]\, Y => sEmpty_RNO_6_2);
    
    \Raddr_vect_RNIQU6A4[4]\ : OA1A
      port map(A => data_mem_ren_i_0(1), B => 
        \data_mem_addr_r_1[4]\, C => N_43, Y => 
        \data_addr_r_iv_i_4[4]\);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_9_0, B => \data_mem_addr_r_1[3]\, Y => 
        I_13_18);
    
    un26_sfull_s_tz_RNO_1 : XA1B
      port map(A => \data_mem_addr_r_1[0]\, B => 
        \un8_waddr_vect_s[0]\, C => data_wen(1), Y => 
        un5_sfull_s_4_0);
    
    \ready_gen.un69_ready_0_I_10\ : OA1A
      port map(A => N_8, B => N_10, C => N_9_1, Y => N_13_0);
    
    \ready_gen.un69_ready_0_I_11\ : OA1
      port map(A => N_13_0, B => N_12_2, C => N_11, Y => 
        un69_ready);
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => \data_mem_addr_w_1[2]\, S
         => data_mem_wen_i_0(1), Y => Waddr_vect_e2);
    
    un60_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0_0 : AO1C
      port map(A => \data_mem_addr_r_1[2]\, B => 
        \data_mem_addr_w_1[2]\, C => N_109, Y => 
        ADD_5x5_fast_I11_Y_i_a2_0);
    
    \Waddr_vect_RNIBOBV[0]\ : OR3A
      port map(A => N_165, B => data_mem_wen_i_0(1), C => 
        \data_mem_addr_w_1[0]\, Y => N_158);
    
    sEmpty_RNO_2 : NOR3C
      port map(A => un7_sempty_s_1, B => un7_sempty_s_0, C => 
        un7_sempty_s_2, Y => un7_sempty_s_4);
    
    un60_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3 : NOR2A
      port map(A => N_9, B => \data_mem_addr_r_1[2]\, Y => N_17);
    
    sEmpty_RNO_4 : XA1A
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \un10_raddr_vect_s[0]\, C => data_wen(1), Y => 
        un7_sempty_s_0);
    
    un75_ready_1_16_ADD_5x5_fast_I11_un1_Y : AOI1B
      port map(A => N_109, B => N_89_i, C => 
        ADD_5x5_fast_I11_un1_Y_0, Y => I11_un1_Y);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_r_1[0]\, B => 
        \data_mem_addr_r_1[1]\, Y => I_5_18);
    
    \Raddr_vect_RNITJRC[4]\ : NOR2B
      port map(A => I_9_18, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[2]\);
    
    \ready_gen.un69_ready_0_I_6\ : OA1A
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \data_mem_addr_r_1[3]\, C => N_5, Y => N_9_1);
    
    un26_sfull_s_tz_RNO_2 : XA1
      port map(A => \data_mem_addr_r_1[3]\, B => 
        \un8_waddr_vect_s[3]\, C => \un26_sfull_s_tz_RNO_7\, Y
         => un5_sfull_s_4_2);
    
    un60_ready_1_1_0_CO1_tz : AO18
      port map(A => N_105_1, B => \data_mem_addr_w_1[2]\, C => 
        \data_mem_addr_r_1[2]\, Y => CO1_tz);
    
    \ready_gen.un69_ready_0_I_3\ : NOR2A
      port map(A => \data_mem_addr_r_1[0]\, B => 
        \data_mem_addr_w_1[0]\, Y => N_6);
    
    sEmpty : DFN1P0
      port map(D => sEmpty_RNO_11, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \sEmpty\);
    
    \Raddr_vect_RNIRSIG2[0]\ : MX2C
      port map(A => \un75_ready1[5]\, B => N_16_i_i_0, S => 
        \data_mem_addr_r_1[0]\, Y => N_197);
    
    \Raddr_vect_RNI4A0PH[0]\ : NOR3C
      port map(A => \data_addr_r_iv_i_4[0]\, B => 
        data_addr_r_iv_i_3(0), C => N_76, Y => 
        Raddr_vect_RNI4A0PH(0));
    
    un75_ready_1_16_ADD_5x5_fast_I16_Y_0 : AX1D
      port map(A => I11_un1_Y, B => ADD_5x5_fast_I11_Y_0, C => 
        N_75_i_0, Y => \un75_ready1[5]\);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \data_mem_addr_w_1[1]\, 
        S => data_mem_wen_i_0(1), Y => Waddr_vect_e1);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_1[2]\);
    
    un6_waddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \data_mem_addr_w_1[1]\, C => \data_mem_addr_w_1[2]\, Y
         => \DWACT_FINC_E[0]\);
    
    \Raddr_vect_RNI7873_0[3]\ : OR2A
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \data_mem_addr_r_1[3]\, Y => N_109);
    
    \Raddr_vect_RNI1473[3]\ : NOR2
      port map(A => \data_mem_addr_r_1[3]\, B => 
        \data_mem_addr_r_1[2]\, Y => un2_raddr_vect_slto3_0);
    
    \Raddr_vect[3]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => data_mem_ren_i_0(1), Q => 
        \data_mem_addr_r_1[3]\);
    
    \Raddr_vect_RNIIMQ5I[4]\ : NOR3C
      port map(A => \data_addr_r_iv_i_4[4]\, B => 
        data_addr_r_iv_i_3(4), C => N_44, Y => 
        Raddr_vect_RNIIMQ5I(4));
    
    sEmpty_RNO_5 : XA1A
      port map(A => \data_mem_addr_w_1[3]\, B => 
        \un10_raddr_vect_s[3]\, C => sEmpty_RNO_7_0, Y => 
        un7_sempty_s_2);
    
    un75_ready_1_16_ADD_5x5_fast_I1_G0N : AO1C
      port map(A => \data_mem_addr_w_1[2]\, B => 
        \data_mem_addr_r_1[2]\, C => N_87, Y => N80);
    
    un8_raddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_r_1[3]\, B => 
        \DWACT_FINC_E_0[0]\, Y => N_4_0);
    
    un60_ready_0_0_0_ADD_5x5_fast_I18_Y_0 : AX1C
      port map(A => N_12_1, B => N_13, C => N_89_i, Y => 
        \un60_ready0[4]\);
    
    un75_ready_1_16_ADD_5x5_fast_I15_Y_0 : AX1A
      port map(A => ADD_5x5_fast_I8_un1_Y_0, B => N80, C => 
        \un75_ready0_1[4]\, Y => \un75_ready1[4]\);
    
    \Raddr_vect[4]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => data_mem_ren_i_0(1), Q => 
        \data_mem_addr_r_1[4]\);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_12, B => \data_mem_addr_w_1[2]\, Y => 
        I_9_17);
    
    un75_ready_1_16_ADD_5x5_fast_I11_Y_0 : MIN3
      port map(A => N_89_i, B => N_109, C => N80, Y => 
        ADD_5x5_fast_I11_Y_0);
    
    sEmpty_RNO_1 : NOR2B
      port map(A => \sEmpty\, B => data_wen(1), Y => un1_sempty_s);
    
    sFull_RNICGOT : OR3B
      port map(A => data_mem_wen_i_0(1), B => data_mem_wen_i_0(2), 
        C => N_164, Y => N_120_i);
    
    \Waddr_vect_RNO_1[2]\ : AX1C
      port map(A => \data_mem_addr_w_1[0]\, B => 
        \data_mem_addr_w_1[1]\, C => \data_mem_addr_w_1[2]\, Y
         => Waddr_vect_n2_tz);
    
    \Raddr_vect_RNIME6A4[2]\ : OA1A
      port map(A => data_mem_ren_i_0(1), B => 
        \data_mem_addr_r_1[2]\, C => N_59, Y => 
        \data_addr_r_iv_i_4[2]\);
    
    un8_raddr_vect_s_I_20 : XOR2
      port map(A => N_4_0, B => \data_mem_addr_r_1[4]\, Y => 
        I_20_10);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ7 is

    port( time_mem_addr_w_3_i_0_1     : out   std_logic;
          data_addr_w_1_iv_i_a2_1_1_0 : in    std_logic_vector(6 to 6);
          data_addr_w_1_iv_i_s_0_0    : out   std_logic_vector(6 to 6);
          time_wen                    : in    std_logic_vector(3 to 3);
          time_ren                    : in    std_logic_vector(3 to 3);
          data_mem_ren_i_0            : in    std_logic_vector(1 to 1);
          time_mem_ren_i_0            : out   std_logic_vector(3 to 3);
          data_addr_r_1_iv_i_a9_1_1   : out   std_logic_vector(6 to 6);
          time_mem_addr_w_3           : out   std_logic_vector(1 downto 0);
          HRESETn_c                   : in    std_logic;
          HCLK_c                      : in    std_logic;
          N_124                       : out   std_logic;
          N_64                        : out   std_logic;
          N_140                       : out   std_logic;
          N_30_1                      : out   std_logic;
          N_89                        : out   std_logic;
          N_163                       : in    std_logic;
          N_164                       : out   std_logic;
          N_72                        : out   std_logic;
          N_56                        : out   std_logic;
          N_48                        : out   std_logic;
          N_35                        : out   std_logic;
          N_113                       : in    std_logic;
          N_162                       : in    std_logic;
          N_77                        : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ7;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ7 is 

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_7, \time_mem_addr_r_3[1]\, \time_mem_addr_r_3[0]\, 
        N_7_0, un5_sfull_s_3, sFull_RNO_3_0, sFull_RNO_4_0, 
        un5_sfull_s_0, un5_sfull_s_2, \Raddr_vect[3]_net_1\, 
        \un8_waddr_vect_s[3]\, \un8_waddr_vect_s[0]\, 
        un7_sempty_s_3, sEmpty_RNO_3_2, sEmpty_RNO_4_2, 
        un7_sempty_s_0, un7_sempty_s_2, \Waddr_vect[3]_net_1\, 
        \un10_raddr_vect_s[3]\, \un10_raddr_vect_s[0]\, 
        \time_mem_addr_w_3[0]\, \data_addr_w_1_iv_i_s_0_tz[6]\, 
        un2_raddr_vect_slt3, \time_mem_addr_r_3_i_0[2]\, 
        un1_waddr_vect_slt3, \time_mem_addr_w_3[1]\, 
        \time_mem_addr_w_3_i_0[2]\, Raddr_vect_n3, Raddr_vect_7_0, 
        Waddr_vect_n3, Waddr_vect_15_0, 
        \time_mem_addr_w_3_i_0[5]\, \time_mem_wen_i_0[3]\, 
        Raddr_vect_n2, un2_raddr_vect_s, Raddr_vect_n2_tz, 
        Waddr_vect_n2, un1_waddr_vect_s, Waddr_vect_n2_tz, I_13_3, 
        I_5_3, I_9_3, \time_mem_addr_r_3_i_0[5]\, 
        \time_mem_ren_i_0[3]\, \time_mem_addr_r_3_i_0[3]\, 
        Raddr_vect_n1_i, Raddr_vect_e2, Raddr_vect_e1, 
        Raddr_vect_e0, \N_89\, Waddr_vect_e2, Waddr_vect_e0, 
        Waddr_vect_e1, Waddr_vect_n1_i, I_13_4, I_5_4, I_9_4, 
        \sFull_RNO\, un8_sfull_s, \sEmpty_RNO\, un2_sempty_s, 
        \sFull\, \sEmpty\, N_4, N_4_0, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    time_mem_ren_i_0(3) <= \time_mem_ren_i_0[3]\;
    time_mem_addr_w_3(1) <= \time_mem_addr_w_3[1]\;
    time_mem_addr_w_3(0) <= \time_mem_addr_w_3[0]\;
    N_89 <= \N_89\;

    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_w_3[1]\, B => 
        \time_mem_addr_w_3[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_w_3[0]\, B => 
        \time_mem_addr_w_3[1]\, C => \time_mem_addr_w_3_i_0[2]\, 
        Y => N_4);
    
    \Raddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_r_3[1]\, B => 
        \time_mem_addr_r_3[0]\, C => un2_raddr_vect_s, Y => 
        Raddr_vect_n1_i);
    
    \Raddr_vect_RNICJ9L[2]\ : OR2A
      port map(A => \time_mem_addr_r_3_i_0[2]\, B => 
        \time_mem_ren_i_0[3]\, Y => N_56);
    
    sFull_RNIR3CG : OR2B
      port map(A => \time_mem_addr_w_3_i_0[5]\, B => \N_89\, Y
         => N_124);
    
    sEmpty_RNIBEFO_1 : OR2
      port map(A => \time_mem_ren_i_0[3]\, B => 
        \time_mem_addr_r_3_i_0[5]\, Y => N_30_1);
    
    \Waddr_vect_RNI6PG9[1]\ : OR3
      port map(A => \time_mem_addr_w_3[0]\, B => 
        \time_mem_addr_w_3[1]\, C => \time_mem_addr_w_3_i_0[2]\, 
        Y => un1_waddr_vect_slt3);
    
    un43_mem_addr_ren_1_SUM1_0 : XNOR2
      port map(A => \time_mem_addr_r_3_i_0[2]\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_3_i_0[3]\);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_w_3[1]\, B => 
        \time_mem_addr_w_3[0]\, Y => N_7_0);
    
    sEmpty_RNO : AO1
      port map(A => un7_sempty_s_3, B => un7_sempty_s_2, C => 
        un2_sempty_s, Y => \sEmpty_RNO\);
    
    \Raddr_vect[1]\ : DFN1C0
      port map(D => Raddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_3[1]\);
    
    \Waddr_vect[3]\ : DFN1E0C0
      port map(D => Waddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_wen_i_0[3]\, Q => 
        \Waddr_vect[3]_net_1\);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_7, B => \time_mem_addr_r_3_i_0[2]\, Y => 
        I_9_4);
    
    sEmpty : DFN1P0
      port map(D => \sEmpty_RNO\, CLK => HCLK_c, PRE => HRESETn_c, 
        Q => \sEmpty\);
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => \time_mem_wen_i_0[3]\, 
        C => \time_mem_addr_w_3[0]\, Y => Waddr_vect_e0);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_3_i_0[2]\);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \time_mem_addr_w_3[1]\, 
        S => \time_mem_wen_i_0[3]\, Y => Waddr_vect_e1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Waddr_vect_RNO_0[2]\ : OR2B
      port map(A => un1_waddr_vect_s, B => Waddr_vect_n2_tz, Y
         => Waddr_vect_n2);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_w_3[0]\, B => 
        \time_mem_addr_w_3[1]\, Y => I_5_3);
    
    \Raddr_vect_RNIMJMC[3]\ : OR2B
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, Y => un2_raddr_vect_s);
    
    \Raddr_vect_RNO_0[2]\ : OR2B
      port map(A => un2_raddr_vect_s, B => Raddr_vect_n2_tz, Y
         => Raddr_vect_n2);
    
    sEmpty_RNIFCRP3 : NOR3B
      port map(A => N_77, B => \time_mem_ren_i_0[3]\, C => 
        data_mem_ren_i_0(1), Y => data_addr_r_1_iv_i_a9_1_1(6));
    
    \Waddr_vect_RNIN86D[2]\ : OR2B
      port map(A => \time_mem_addr_w_3_i_0[2]\, B => \N_89\, Y
         => N_140);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => Raddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_ren_i_0[3]\, Q => 
        \Raddr_vect[3]_net_1\);
    
    sEmpty_RNO_2 : NOR2B
      port map(A => time_wen(3), B => \sEmpty\, Y => un2_sempty_s);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_4, B => \Waddr_vect[3]_net_1\, Y => I_13_3);
    
    sFull_RNO : AO1
      port map(A => un5_sfull_s_3, B => un5_sfull_s_2, C => 
        un8_sfull_s, Y => \sFull_RNO\);
    
    \Raddr_vect_RNO[0]\ : AXOI7
      port map(A => un2_raddr_vect_s, B => \time_mem_ren_i_0[3]\, 
        C => \time_mem_addr_r_3[0]\, Y => Raddr_vect_e0);
    
    \Raddr_vect_RNO[1]\ : MX2A
      port map(A => Raddr_vect_n1_i, B => \time_mem_addr_r_3[1]\, 
        S => \time_mem_ren_i_0[3]\, Y => Raddr_vect_e1);
    
    sFull_RNIKH0A_0 : NOR2A
      port map(A => N_163, B => \time_mem_wen_i_0[3]\, Y => 
        \N_89\);
    
    sFull_RNO_4 : AX1E
      port map(A => un1_waddr_vect_s, B => I_5_3, C => 
        \time_mem_addr_r_3[1]\, Y => sFull_RNO_4_0);
    
    sFull_RNO_6 : OR2B
      port map(A => I_13_3, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    sEmpty_RNO_3 : AX1E
      port map(A => un2_raddr_vect_s, B => I_9_4, C => 
        \time_mem_addr_w_3_i_0[2]\, Y => sEmpty_RNO_3_2);
    
    \Raddr_vect[2]\ : DFN1C0
      port map(D => Raddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_3_i_0[2]\);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_3[0]\);
    
    sFull_RNO_5 : XA1B
      port map(A => \un8_waddr_vect_s[0]\, B => 
        \time_mem_addr_r_3[0]\, C => time_wen(3), Y => 
        un5_sfull_s_0);
    
    sFull_RNIQOVC1 : OA1
      port map(A => N_162, B => \data_addr_w_1_iv_i_s_0_tz[6]\, C
         => N_113, Y => data_addr_w_1_iv_i_s_0_0(6));
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => 
        \time_mem_addr_w_3_i_0[2]\, S => \time_mem_wen_i_0[3]\, Y
         => Waddr_vect_e2);
    
    sEmpty_RNO_4 : AX1E
      port map(A => un2_raddr_vect_s, B => I_5_4, C => 
        \time_mem_addr_w_3[1]\, Y => sEmpty_RNO_4_2);
    
    un50_mem_addr_wen_1_SUM1_0 : XNOR2
      port map(A => \time_mem_addr_w_3_i_0[2]\, B => 
        \Waddr_vect[3]_net_1\, Y => time_mem_addr_w_3_i_0_1);
    
    sFull_RNO_3 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_3, C => 
        \time_mem_addr_r_3_i_0[2]\, Y => sFull_RNO_3_0);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => sEmpty_RNO_3_2, B => sEmpty_RNO_4_2, C => 
        un7_sempty_s_0, Y => un7_sempty_s_3);
    
    \Waddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_w_3[0]\, B => 
        \time_mem_addr_w_3[1]\, C => \time_mem_addr_w_3_i_0[2]\, 
        Y => Waddr_vect_n2_tz);
    
    \Raddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_r_3[0]\, B => 
        \time_mem_addr_r_3[1]\, C => \time_mem_addr_r_3_i_0[2]\, 
        Y => Raddr_vect_n2_tz);
    
    sEmpty_RNO_7 : OR2A
      port map(A => un2_raddr_vect_s, B => \time_mem_addr_r_3[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Raddr_vect_RNO[2]\ : MX2A
      port map(A => Raddr_vect_n2, B => 
        \time_mem_addr_r_3_i_0[2]\, S => \time_mem_ren_i_0[3]\, Y
         => Raddr_vect_e2);
    
    \Raddr_vect[0]\ : DFN1C0
      port map(D => Raddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_3[0]\);
    
    sEmpty_RNIBEFO_0 : OR2A
      port map(A => \time_mem_addr_r_3_i_0[3]\, B => 
        \time_mem_ren_i_0[3]\, Y => N_48);
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_r_3[1]\, B => 
        \time_mem_addr_r_3[0]\, Y => N_7);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_7_0, B => \time_mem_addr_w_3_i_0[2]\, Y => 
        I_9_3);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_4_0, B => \Raddr_vect[3]_net_1\, Y => 
        I_13_4);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_r_3[0]\, B => 
        \time_mem_addr_r_3[1]\, C => \time_mem_addr_r_3_i_0[2]\, 
        Y => N_4_0);
    
    sFull_RNIBLJS : MX2B
      port map(A => \time_mem_addr_w_3_i_0[5]\, B => 
        data_addr_w_1_iv_i_a2_1_1_0(6), S => 
        \time_mem_wen_i_0[3]\, Y => 
        \data_addr_w_1_iv_i_s_0_tz[6]\);
    
    sFull_RNIG4G2 : OR2
      port map(A => time_wen(3), B => \sFull\, Y => 
        \time_mem_wen_i_0[3]\);
    
    \Raddr_vect_RNINOG9[1]\ : OR3
      port map(A => \time_mem_addr_r_3[0]\, B => 
        \time_mem_addr_r_3[1]\, C => \time_mem_addr_r_3_i_0[2]\, 
        Y => un2_raddr_vect_slt3);
    
    sEmpty_RNO_1 : XA1B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \un10_raddr_vect_s[3]\, C => time_ren(3), Y => 
        un7_sempty_s_2);
    
    sFull_RNO_1 : XA1
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \un8_waddr_vect_s[3]\, C => time_ren(3), Y => 
        un5_sfull_s_2);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_r_3[0]\, B => 
        \time_mem_addr_r_3[1]\, Y => I_5_4);
    
    \Waddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_w_3[0]\, B => 
        \time_mem_addr_w_3[1]\, C => \time_mem_addr_w_3_i_0[2]\, 
        Y => Waddr_vect_15_0);
    
    sFull_RNO_7 : OR2A
      port map(A => un1_waddr_vect_s, B => \time_mem_addr_w_3[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    sEmpty_RNIBEFO : OR2A
      port map(A => \time_mem_addr_r_3_i_0[5]\, B => 
        \time_mem_ren_i_0[3]\, Y => N_35);
    
    \Raddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_r_3[0]\, B => 
        \time_mem_addr_r_3[1]\, C => \time_mem_addr_r_3_i_0[2]\, 
        Y => Raddr_vect_7_0);
    
    \Waddr_vect_RNO[3]\ : AXOI1
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, C => Waddr_vect_15_0, Y => 
        Waddr_vect_n3);
    
    sFull_RNO_0 : NOR3C
      port map(A => sFull_RNO_3_0, B => sFull_RNO_4_0, C => 
        un5_sfull_s_0, Y => un5_sfull_s_3);
    
    sEmpty_RNO_6 : OR2B
      port map(A => I_13_4, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    un43_mem_addr_ren_1_CO1 : NOR2B
      port map(A => \time_mem_addr_r_3_i_0[2]\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_3_i_0[5]\);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => \sFull\);
    
    \Waddr_vect_RNIAKMC[3]\ : OR2B
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, Y => un1_waddr_vect_s);
    
    un50_mem_addr_wen_1_CO1 : NOR2B
      port map(A => \time_mem_addr_w_3_i_0[2]\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_3_i_0[5]\);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_3[1]\);
    
    sEmpty_RNIES3I : OR2
      port map(A => time_ren(3), B => \sEmpty\, Y => 
        \time_mem_ren_i_0[3]\);
    
    \Raddr_vect_RNIBF9L[1]\ : OR2
      port map(A => \time_mem_ren_i_0[3]\, B => 
        \time_mem_addr_r_3[1]\, Y => N_64);
    
    sFull_RNO_2 : NOR2B
      port map(A => time_ren(3), B => \sFull\, Y => un8_sfull_s);
    
    sEmpty_RNO_5 : XA1
      port map(A => \un10_raddr_vect_s[0]\, B => 
        \time_mem_addr_w_3[0]\, C => time_wen(3), Y => 
        un7_sempty_s_0);
    
    \Raddr_vect_RNO[3]\ : AXOI1
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, C => Raddr_vect_7_0, Y => 
        Raddr_vect_n3);
    
    \Raddr_vect_RNIAB9L[0]\ : OR2
      port map(A => \time_mem_ren_i_0[3]\, B => 
        \time_mem_addr_r_3[0]\, Y => N_72);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    sFull_RNIKH0A : OR2B
      port map(A => \time_mem_wen_i_0[3]\, B => N_163, Y => N_164);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity generic_syncram_2p_7_32_0 is

    port( wdata                         : in    std_logic_vector(31 downto 0);
          Waddr_vect_RNILLSP5           : in    std_logic_vector(4 to 4);
          Waddr_vect_RNIJTNE5           : in    std_logic_vector(3 to 3);
          Waddr_vect_RNI394D5           : in    std_logic_vector(2 to 2);
          Waddr_vect_RNI0O455           : in    std_logic_vector(1 to 1);
          Waddr_vect_RNION355           : in    std_logic_vector(0 to 0);
          Raddr_vect_RNIIMQ5I           : in    std_logic_vector(4 to 4);
          Raddr_vect_RNIE6Q5I           : in    std_logic_vector(3 to 3);
          Raddr_vect_RNIKA2PH           : in    std_logic_vector(2 to 2);
          Raddr_vect_RNICA1PH           : in    std_logic_vector(1 to 1);
          Raddr_vect_RNI4A0PH           : in    std_logic_vector(0 to 0);
          hwdata_c                      : out   std_logic_vector(31 downto 0);
          N_1_i_1_i                     : in    std_logic;
          generic_syncram_2p_7_32_0_VCC : in    std_logic;
          generic_syncram_2p_7_32_0_GND : in    std_logic;
          sFull_RNIU5GK1                : in    std_logic;
          sFull_RNIHL443                : in    std_logic;
          sEmpty_RNILSD08               : in    std_logic;
          sEmpty_RNIE7T87               : in    std_logic;
          N_1_i_1                       : in    std_logic;
          HCLK_c                        : in    std_logic
        );

end generic_syncram_2p_7_32_0;

architecture DEF_ARCH of generic_syncram_2p_7_32_0 is 

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM512X18
    generic (MEMORYFILE:string := "");

    port( RADDR8 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          WADDR8 : in    std_logic := 'U';
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          WD17   : in    std_logic := 'U';
          WD16   : in    std_logic := 'U';
          WD15   : in    std_logic := 'U';
          WD14   : in    std_logic := 'U';
          WD13   : in    std_logic := 'U';
          WD12   : in    std_logic := 'U';
          WD11   : in    std_logic := 'U';
          WD10   : in    std_logic := 'U';
          WD9    : in    std_logic := 'U';
          WD8    : in    std_logic := 'U';
          WD7    : in    std_logic := 'U';
          WD6    : in    std_logic := 'U';
          WD5    : in    std_logic := 'U';
          WD4    : in    std_logic := 'U';
          WD3    : in    std_logic := 'U';
          WD2    : in    std_logic := 'U';
          WD1    : in    std_logic := 'U';
          WD0    : in    std_logic := 'U';
          RW0    : in    std_logic := 'U';
          RW1    : in    std_logic := 'U';
          WW0    : in    std_logic := 'U';
          WW1    : in    std_logic := 'U';
          PIPE   : in    std_logic := 'U';
          REN    : in    std_logic := 'U';
          WEN    : in    std_logic := 'U';
          RCLK   : in    std_logic := 'U';
          WCLK   : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          RD17   : out   std_logic;
          RD16   : out   std_logic;
          RD15   : out   std_logic;
          RD14   : out   std_logic;
          RD13   : out   std_logic;
          RD12   : out   std_logic;
          RD11   : out   std_logic;
          RD10   : out   std_logic;
          RD9    : out   std_logic;
          RD8    : out   std_logic;
          RD7    : out   std_logic;
          RD6    : out   std_logic;
          RD5    : out   std_logic;
          RD4    : out   std_logic;
          RD3    : out   std_logic;
          RD2    : out   std_logic;
          RD1    : out   std_logic;
          RD0    : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_7_0, I_5_1, I_5_0, I_5_5, I_4_5_i_0, I_4_4_i_0, 
        I_5_3, \RADDR_REG1[6]\, \WADDR_REG1[6]\, N_5, 
        \RADDR_REG1[2]\, \WADDR_REG1[2]\, I_4_3_i_0, 
        \RADDR_REG1[0]\, \WADDR_REG1[0]\, I_4_1_i_0, N_7, 
        \DOUT_TMP[13]\, \DIN_REG1[13]\, \DOUT_TMP[12]\, 
        \DIN_REG1[12]\, \DOUT_TMP[11]\, \DIN_REG1[11]\, 
        \DOUT_TMP[10]\, \DIN_REG1[10]\, \DOUT_TMP[9]\, 
        \DIN_REG1[9]\, \DOUT_TMP[8]\, \DIN_REG1[8]\, 
        \DOUT_TMP[7]\, \DIN_REG1[7]\, \DOUT_TMP[6]\, 
        \DIN_REG1[6]\, \DOUT_TMP[5]\, \DIN_REG1[5]\, 
        \DOUT_TMP[4]\, \DIN_REG1[4]\, \DOUT_TMP[3]\, 
        \DIN_REG1[3]\, \DOUT_TMP[2]\, \DIN_REG1[2]\, 
        \DOUT_TMP[1]\, \DIN_REG1[1]\, \DOUT_TMP[0]\, 
        \DIN_REG1[0]\, \DOUT_TMP[17]\, \DIN_REG1[17]\, 
        \DOUT_TMP[16]\, \DIN_REG1[16]\, \DOUT_TMP[15]\, 
        \DIN_REG1[15]\, \DOUT_TMP[14]\, \DIN_REG1[14]\, 
        \DOUT_TMP_0[13]\, \DIN_REG1_0[13]\, \DOUT_TMP_0[12]\, 
        \DIN_REG1_0[12]\, \DOUT_TMP_0[11]\, \DIN_REG1_0[11]\, 
        \DOUT_TMP_0[10]\, \DIN_REG1_0[10]\, \DOUT_TMP_0[9]\, 
        \DIN_REG1_0[9]\, \DOUT_TMP_0[8]\, \DIN_REG1_0[8]\, 
        \DOUT_TMP_0[7]\, \DIN_REG1_0[7]\, \DOUT_TMP_0[6]\, 
        \DIN_REG1_0[6]\, \DOUT_TMP_0[5]\, \DIN_REG1_0[5]\, 
        \DOUT_TMP_0[4]\, \DIN_REG1_0[4]\, \DOUT_TMP_0[3]\, 
        \DIN_REG1_0[3]\, \DOUT_TMP_0[2]\, \DIN_REG1_0[2]\, 
        \DOUT_TMP_0[1]\, \DIN_REG1_0[1]\, \DOUT_TMP_0[0]\, 
        \DIN_REG1_0[0]\, \WADDR_REG1[5]\, \RADDR_REG1[5]\, 
        \WADDR_REG1[4]\, \RADDR_REG1[4]\, \WADDR_REG1[3]\, 
        \RADDR_REG1[3]\, \WADDR_REG1[1]\, \RADDR_REG1[1]\, 
        \DOUT_TMP_0[14]\, \DOUT_TMP_0[15]\, \DOUT_TMP_0[16]\, 
        \DOUT_TMP_0[17]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \rfd_tile_RADDR_REG1_RNIG9I4[2]\ : XA1A
      port map(A => \RADDR_REG1[2]\, B => \WADDR_REG1[2]\, C => 
        I_4_3_i_0, Y => I_5_1);
    
    \rfd_tile_DIN_REG1[9]\ : DFN1
      port map(D => wdata(9), CLK => HCLK_c, Q => \DIN_REG1_0[9]\);
    
    \rfd_tile_0_DIN_REG1[0]\ : DFN1
      port map(D => wdata(18), CLK => HCLK_c, Q => \DIN_REG1[0]\);
    
    \rfd_tile_RADDR_REG1[5]\ : DFN1
      port map(D => sEmpty_RNIE7T87, CLK => HCLK_c, Q => 
        \RADDR_REG1[5]\);
    
    \rfd_tile_0_DIN_REG1[12]\ : DFN1
      port map(D => wdata(30), CLK => HCLK_c, Q => \DIN_REG1[12]\);
    
    \rfd_tile_WADDR_REG1[6]\ : DFN1
      port map(D => sFull_RNIU5GK1, CLK => HCLK_c, Q => 
        \WADDR_REG1[6]\);
    
    rfd_tile_I_3 : DFN1
      port map(D => N_1_i_1, CLK => HCLK_c, Q => N_5);
    
    \rfd_tile_RADDR_REG1_RNI89H4[0]\ : XA1A
      port map(A => \RADDR_REG1[0]\, B => \WADDR_REG1[0]\, C => 
        I_4_1_i_0, Y => I_5_0);
    
    rfd_tile_0_I_1_RNIK6BO : MX2
      port map(A => \DOUT_TMP[6]\, B => \DIN_REG1[6]\, S => N_7_0, 
        Y => hwdata_c(24));
    
    rfd_tile_I_1_RNI83001 : MX2
      port map(A => \DOUT_TMP_0[13]\, B => \DIN_REG1_0[13]\, S
         => N_7, Y => hwdata_c(13));
    
    \rfd_tile_0_DIN_REG1[11]\ : DFN1
      port map(D => wdata(29), CLK => HCLK_c, Q => \DIN_REG1[11]\);
    
    \rfd_tile_DIN_REG1[10]\ : DFN1
      port map(D => wdata(10), CLK => HCLK_c, Q => 
        \DIN_REG1_0[10]\);
    
    rfd_tile_0_I_1_RNIGMAO : MX2
      port map(A => \DOUT_TMP[2]\, B => \DIN_REG1[2]\, S => N_7_0, 
        Y => hwdata_c(20));
    
    rfd_tile_I_1_RNIA3001 : MX2
      port map(A => \DOUT_TMP[15]\, B => \DIN_REG1[15]\, S => N_7, 
        Y => hwdata_c(15));
    
    \rfd_tile_DIN_REG1_RNIROBR[7]\ : MX2
      port map(A => \DOUT_TMP_0[7]\, B => \DIN_REG1_0[7]\, S => 
        N_7, Y => hwdata_c(7));
    
    \rfd_tile_WADDR_REG1[4]\ : DFN1
      port map(D => Waddr_vect_RNILLSP5(4), CLK => HCLK_c, Q => 
        \WADDR_REG1[4]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \rfd_tile_DIN_REG1_RNIM4BR[2]\ : MX2
      port map(A => \DOUT_TMP_0[2]\, B => \DIN_REG1_0[2]\, S => 
        N_7, Y => hwdata_c(2));
    
    \rfd_tile_DIN_REG1[0]\ : DFN1
      port map(D => wdata(0), CLK => HCLK_c, Q => \DIN_REG1_0[0]\);
    
    \rfd_tile_DIN_REG1[5]\ : DFN1
      port map(D => wdata(5), CLK => HCLK_c, Q => \DIN_REG1_0[5]\);
    
    \rfd_tile_0_DIN_REG1[6]\ : DFN1
      port map(D => wdata(24), CLK => HCLK_c, Q => \DIN_REG1[6]\);
    
    \rfd_tile_0_DIN_REG1[1]\ : DFN1
      port map(D => wdata(19), CLK => HCLK_c, Q => \DIN_REG1[1]\);
    
    \rfd_tile_RADDR_REG1_RNILO82[1]\ : XNOR2
      port map(A => \WADDR_REG1[1]\, B => \RADDR_REG1[1]\, Y => 
        I_4_1_i_0);
    
    \rfd_tile_DIN_REG1[4]\ : DFN1
      port map(D => wdata(4), CLK => HCLK_c, Q => \DIN_REG1_0[4]\);
    
    \rfd_tile_DIN_REG1[3]\ : DFN1
      port map(D => wdata(3), CLK => HCLK_c, Q => \DIN_REG1_0[3]\);
    
    \rfd_tile_DIN_REG1[2]\ : DFN1
      port map(D => wdata(2), CLK => HCLK_c, Q => \DIN_REG1_0[2]\);
    
    rfd_tile_0_I_1_RNIHQAO : MX2
      port map(A => \DOUT_TMP[3]\, B => \DIN_REG1[3]\, S => N_7_0, 
        Y => hwdata_c(21));
    
    \rfd_tile_0_DIN_REG1[2]\ : DFN1
      port map(D => wdata(20), CLK => HCLK_c, Q => \DIN_REG1[2]\);
    
    rfd_tile_0_I_1 : RAM512X18
      port map(RADDR8 => generic_syncram_2p_7_32_0_GND, RADDR7
         => generic_syncram_2p_7_32_0_GND, RADDR6 => 
        sEmpty_RNILSD08, RADDR5 => sEmpty_RNIE7T87, RADDR4 => 
        Raddr_vect_RNIIMQ5I(4), RADDR3 => Raddr_vect_RNIE6Q5I(3), 
        RADDR2 => Raddr_vect_RNIKA2PH(2), RADDR1 => 
        Raddr_vect_RNICA1PH(1), RADDR0 => Raddr_vect_RNI4A0PH(0), 
        WADDR8 => generic_syncram_2p_7_32_0_GND, WADDR7 => 
        generic_syncram_2p_7_32_0_GND, WADDR6 => sFull_RNIU5GK1, 
        WADDR5 => sFull_RNIHL443, WADDR4 => 
        Waddr_vect_RNILLSP5(4), WADDR3 => Waddr_vect_RNIJTNE5(3), 
        WADDR2 => Waddr_vect_RNI394D5(2), WADDR1 => 
        Waddr_vect_RNI0O455(1), WADDR0 => Waddr_vect_RNION355(0), 
        WD17 => generic_syncram_2p_7_32_0_GND, WD16 => 
        generic_syncram_2p_7_32_0_GND, WD15 => 
        generic_syncram_2p_7_32_0_GND, WD14 => 
        generic_syncram_2p_7_32_0_GND, WD13 => wdata(31), WD12
         => wdata(30), WD11 => wdata(29), WD10 => wdata(28), WD9
         => wdata(27), WD8 => wdata(26), WD7 => wdata(25), WD6
         => wdata(24), WD5 => wdata(23), WD4 => wdata(22), WD3
         => wdata(21), WD2 => wdata(20), WD1 => wdata(19), WD0
         => wdata(18), RW0 => generic_syncram_2p_7_32_0_GND, RW1
         => generic_syncram_2p_7_32_0_VCC, WW0 => 
        generic_syncram_2p_7_32_0_GND, WW1 => 
        generic_syncram_2p_7_32_0_VCC, PIPE => 
        generic_syncram_2p_7_32_0_GND, REN => 
        generic_syncram_2p_7_32_0_GND, WEN => N_1_i_1_i, RCLK => 
        HCLK_c, WCLK => HCLK_c, RESET => 
        generic_syncram_2p_7_32_0_VCC, RD17 => \DOUT_TMP_0[17]\, 
        RD16 => \DOUT_TMP_0[16]\, RD15 => \DOUT_TMP_0[15]\, RD14
         => \DOUT_TMP_0[14]\, RD13 => \DOUT_TMP[13]\, RD12 => 
        \DOUT_TMP[12]\, RD11 => \DOUT_TMP[11]\, RD10 => 
        \DOUT_TMP[10]\, RD9 => \DOUT_TMP[9]\, RD8 => 
        \DOUT_TMP[8]\, RD7 => \DOUT_TMP[7]\, RD6 => \DOUT_TMP[6]\, 
        RD5 => \DOUT_TMP[5]\, RD4 => \DOUT_TMP[4]\, RD3 => 
        \DOUT_TMP[3]\, RD2 => \DOUT_TMP[2]\, RD1 => \DOUT_TMP[1]\, 
        RD0 => \DOUT_TMP[0]\);
    
    \rfd_tile_DIN_REG1[12]\ : DFN1
      port map(D => wdata(12), CLK => HCLK_c, Q => 
        \DIN_REG1_0[12]\);
    
    \rfd_tile_0_DIN_REG1[5]\ : DFN1
      port map(D => wdata(23), CLK => HCLK_c, Q => \DIN_REG1[5]\);
    
    rfd_tile_0_I_1_RNIMEBO : MX2
      port map(A => \DOUT_TMP[8]\, B => \DIN_REG1[8]\, S => N_7_0, 
        Y => hwdata_c(26));
    
    \rfd_tile_0_DIN_REG1[3]\ : DFN1
      port map(D => wdata(21), CLK => HCLK_c, Q => \DIN_REG1[3]\);
    
    \rfd_tile_RADDR_REG1_RNIRG92[4]\ : XNOR2
      port map(A => \WADDR_REG1[4]\, B => \RADDR_REG1[4]\, Y => 
        I_4_4_i_0);
    
    rfd_tile_0_I_1_RNIIUAO : MX2
      port map(A => \DOUT_TMP[4]\, B => \DIN_REG1[4]\, S => N_7_0, 
        Y => hwdata_c(22));
    
    \rfd_tile_DIN_REG1_RNIPGBR[5]\ : MX2
      port map(A => \DOUT_TMP_0[5]\, B => \DIN_REG1_0[5]\, S => 
        N_7, Y => hwdata_c(5));
    
    rfd_tile_I_1_RNI53001 : MX2
      port map(A => \DOUT_TMP_0[10]\, B => \DIN_REG1_0[10]\, S
         => N_7, Y => hwdata_c(10));
    
    \rfd_tile_DIN_REG1[15]\ : DFN1
      port map(D => wdata(15), CLK => HCLK_c, Q => \DIN_REG1[15]\);
    
    rfd_tile_0_I_1_RNIB01O : MX2
      port map(A => \DOUT_TMP[12]\, B => \DIN_REG1[12]\, S => 
        N_7_0, Y => hwdata_c(30));
    
    \rfd_tile_RADDR_REG1[0]\ : DFN1
      port map(D => Raddr_vect_RNI4A0PH(0), CLK => HCLK_c, Q => 
        \RADDR_REG1[0]\);
    
    \rfd_tile_WADDR_REG1[5]\ : DFN1
      port map(D => sFull_RNIHL443, CLK => HCLK_c, Q => 
        \WADDR_REG1[5]\);
    
    \rfd_tile_RADDR_REG1[2]\ : DFN1
      port map(D => Raddr_vect_RNIKA2PH(2), CLK => HCLK_c, Q => 
        \RADDR_REG1[2]\);
    
    rfd_tile_0_I_1_RNILABO : MX2
      port map(A => \DOUT_TMP[7]\, B => \DIN_REG1[7]\, S => N_7_0, 
        Y => hwdata_c(25));
    
    rfd_tile_0_I_1_RNIFIAO : MX2
      port map(A => \DOUT_TMP[1]\, B => \DIN_REG1[1]\, S => N_7_0, 
        Y => hwdata_c(19));
    
    \rfd_tile_0_DIN_REG1[9]\ : DFN1
      port map(D => wdata(27), CLK => HCLK_c, Q => \DIN_REG1[9]\);
    
    \rfd_tile_DIN_REG1[1]\ : DFN1
      port map(D => wdata(1), CLK => HCLK_c, Q => \DIN_REG1_0[1]\);
    
    \rfd_tile_RADDR_REG1_RNIP892[3]\ : XNOR2
      port map(A => \WADDR_REG1[3]\, B => \RADDR_REG1[3]\, Y => 
        I_4_3_i_0);
    
    rfd_tile_I_1_RNI63001 : MX2
      port map(A => \DOUT_TMP_0[11]\, B => \DIN_REG1_0[11]\, S
         => N_7, Y => hwdata_c(11));
    
    \rfd_tile_RADDR_REG1_RNIQS1L[0]\ : NOR3C
      port map(A => I_5_1, B => I_5_0, C => I_5_5, Y => N_7_0);
    
    \rfd_tile_RADDR_REG1[3]\ : DFN1
      port map(D => Raddr_vect_RNIE6Q5I(3), CLK => HCLK_c, Q => 
        \RADDR_REG1[3]\);
    
    \rfd_tile_DIN_REG1_RNIQKBR[6]\ : MX2
      port map(A => \DOUT_TMP_0[6]\, B => \DIN_REG1_0[6]\, S => 
        N_7, Y => hwdata_c(6));
    
    rfd_tile_0_I_1_RNIJ2BO : MX2
      port map(A => \DOUT_TMP[5]\, B => \DIN_REG1[5]\, S => N_7_0, 
        Y => hwdata_c(23));
    
    \rfd_tile_RADDR_REG1_RNI2AUB[4]\ : NOR3C
      port map(A => I_4_5_i_0, B => I_4_4_i_0, C => I_5_3, Y => 
        I_5_5);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \rfd_tile_RADDR_REG1_RNITO92[5]\ : XNOR2
      port map(A => \WADDR_REG1[5]\, B => \RADDR_REG1[5]\, Y => 
        I_4_5_i_0);
    
    \rfd_tile_RADDR_REG1[1]\ : DFN1
      port map(D => Raddr_vect_RNICA1PH(1), CLK => HCLK_c, Q => 
        \RADDR_REG1[1]\);
    
    \rfd_tile_RADDR_REG1_RNIA0B7[6]\ : XA1A
      port map(A => \RADDR_REG1[6]\, B => \WADDR_REG1[6]\, C => 
        N_5, Y => I_5_3);
    
    rfd_tile_0_I_1_RNINIBO : MX2
      port map(A => \DOUT_TMP[9]\, B => \DIN_REG1[9]\, S => N_7_0, 
        Y => hwdata_c(27));
    
    \rfd_tile_DIN_REG1[14]\ : DFN1
      port map(D => wdata(14), CLK => HCLK_c, Q => \DIN_REG1[14]\);
    
    \rfd_tile_0_DIN_REG1[10]\ : DFN1
      port map(D => wdata(28), CLK => HCLK_c, Q => \DIN_REG1[10]\);
    
    \rfd_tile_DIN_REG1_RNISSBR[8]\ : MX2
      port map(A => \DOUT_TMP_0[8]\, B => \DIN_REG1_0[8]\, S => 
        N_7, Y => hwdata_c(8));
    
    \rfd_tile_RADDR_REG1[6]\ : DFN1
      port map(D => sEmpty_RNILSD08, CLK => HCLK_c, Q => 
        \RADDR_REG1[6]\);
    
    rfd_tile_0_I_1_RNIC01O : MX2
      port map(A => \DOUT_TMP[13]\, B => \DIN_REG1[13]\, S => 
        N_7_0, Y => hwdata_c(31));
    
    rfd_tile_0_I_1_RNIA01O : MX2
      port map(A => \DOUT_TMP[11]\, B => \DIN_REG1[11]\, S => 
        N_7_0, Y => hwdata_c(29));
    
    \rfd_tile_DIN_REG1_RNIKSAR[0]\ : MX2
      port map(A => \DOUT_TMP_0[0]\, B => \DIN_REG1_0[0]\, S => 
        N_7, Y => hwdata_c(0));
    
    \rfd_tile_DIN_REG1_RNIOCBR[4]\ : MX2
      port map(A => \DOUT_TMP_0[4]\, B => \DIN_REG1_0[4]\, S => 
        N_7, Y => hwdata_c(4));
    
    \rfd_tile_DIN_REG1_RNIT0CR[9]\ : MX2
      port map(A => \DOUT_TMP_0[9]\, B => \DIN_REG1_0[9]\, S => 
        N_7, Y => hwdata_c(9));
    
    \rfd_tile_0_DIN_REG1[7]\ : DFN1
      port map(D => wdata(25), CLK => HCLK_c, Q => \DIN_REG1[7]\);
    
    \rfd_tile_0_DIN_REG1[13]\ : DFN1
      port map(D => wdata(31), CLK => HCLK_c, Q => \DIN_REG1[13]\);
    
    \rfd_tile_DIN_REG1[8]\ : DFN1
      port map(D => wdata(8), CLK => HCLK_c, Q => \DIN_REG1_0[8]\);
    
    rfd_tile_0_I_1_RNIEEAO : MX2
      port map(A => \DOUT_TMP[0]\, B => \DIN_REG1[0]\, S => N_7_0, 
        Y => hwdata_c(18));
    
    \rfd_tile_WADDR_REG1[0]\ : DFN1
      port map(D => Waddr_vect_RNION355(0), CLK => HCLK_c, Q => 
        \WADDR_REG1[0]\);
    
    \rfd_tile_DIN_REG1_RNIN8BR[3]\ : MX2
      port map(A => \DOUT_TMP_0[3]\, B => \DIN_REG1_0[3]\, S => 
        N_7, Y => hwdata_c(3));
    
    \rfd_tile_RADDR_REG1[4]\ : DFN1
      port map(D => Raddr_vect_RNIIMQ5I(4), CLK => HCLK_c, Q => 
        \RADDR_REG1[4]\);
    
    \rfd_tile_DIN_REG1[6]\ : DFN1
      port map(D => wdata(6), CLK => HCLK_c, Q => \DIN_REG1_0[6]\);
    
    \rfd_tile_0_DIN_REG1[8]\ : DFN1
      port map(D => wdata(26), CLK => HCLK_c, Q => \DIN_REG1[8]\);
    
    \rfd_tile_WADDR_REG1[2]\ : DFN1
      port map(D => Waddr_vect_RNI394D5(2), CLK => HCLK_c, Q => 
        \WADDR_REG1[2]\);
    
    \rfd_tile_DIN_REG1_RNIL0BR[1]\ : MX2
      port map(A => \DOUT_TMP_0[1]\, B => \DIN_REG1_0[1]\, S => 
        N_7, Y => hwdata_c(1));
    
    \rfd_tile_DIN_REG1[11]\ : DFN1
      port map(D => wdata(11), CLK => HCLK_c, Q => 
        \DIN_REG1_0[11]\);
    
    rfd_tile_I_1_RNI93001 : MX2
      port map(A => \DOUT_TMP[14]\, B => \DIN_REG1[14]\, S => N_7, 
        Y => hwdata_c(14));
    
    \rfd_tile_WADDR_REG1[3]\ : DFN1
      port map(D => Waddr_vect_RNIJTNE5(3), CLK => HCLK_c, Q => 
        \WADDR_REG1[3]\);
    
    \rfd_tile_DIN_REG1[13]\ : DFN1
      port map(D => wdata(13), CLK => HCLK_c, Q => 
        \DIN_REG1_0[13]\);
    
    rfd_tile_0_I_1_RNI901O : MX2
      port map(A => \DOUT_TMP[10]\, B => \DIN_REG1[10]\, S => 
        N_7_0, Y => hwdata_c(28));
    
    rfd_tile_I_1 : RAM512X18
      port map(RADDR8 => generic_syncram_2p_7_32_0_GND, RADDR7
         => generic_syncram_2p_7_32_0_GND, RADDR6 => 
        sEmpty_RNILSD08, RADDR5 => sEmpty_RNIE7T87, RADDR4 => 
        Raddr_vect_RNIIMQ5I(4), RADDR3 => Raddr_vect_RNIE6Q5I(3), 
        RADDR2 => Raddr_vect_RNIKA2PH(2), RADDR1 => 
        Raddr_vect_RNICA1PH(1), RADDR0 => Raddr_vect_RNI4A0PH(0), 
        WADDR8 => generic_syncram_2p_7_32_0_GND, WADDR7 => 
        generic_syncram_2p_7_32_0_GND, WADDR6 => sFull_RNIU5GK1, 
        WADDR5 => sFull_RNIHL443, WADDR4 => 
        Waddr_vect_RNILLSP5(4), WADDR3 => Waddr_vect_RNIJTNE5(3), 
        WADDR2 => Waddr_vect_RNI394D5(2), WADDR1 => 
        Waddr_vect_RNI0O455(1), WADDR0 => Waddr_vect_RNION355(0), 
        WD17 => wdata(17), WD16 => wdata(16), WD15 => wdata(15), 
        WD14 => wdata(14), WD13 => wdata(13), WD12 => wdata(12), 
        WD11 => wdata(11), WD10 => wdata(10), WD9 => wdata(9), 
        WD8 => wdata(8), WD7 => wdata(7), WD6 => wdata(6), WD5
         => wdata(5), WD4 => wdata(4), WD3 => wdata(3), WD2 => 
        wdata(2), WD1 => wdata(1), WD0 => wdata(0), RW0 => 
        generic_syncram_2p_7_32_0_GND, RW1 => 
        generic_syncram_2p_7_32_0_VCC, WW0 => 
        generic_syncram_2p_7_32_0_GND, WW1 => 
        generic_syncram_2p_7_32_0_VCC, PIPE => 
        generic_syncram_2p_7_32_0_GND, REN => 
        generic_syncram_2p_7_32_0_GND, WEN => N_1_i_1_i, RCLK => 
        HCLK_c, WCLK => HCLK_c, RESET => 
        generic_syncram_2p_7_32_0_VCC, RD17 => \DOUT_TMP[17]\, 
        RD16 => \DOUT_TMP[16]\, RD15 => \DOUT_TMP[15]\, RD14 => 
        \DOUT_TMP[14]\, RD13 => \DOUT_TMP_0[13]\, RD12 => 
        \DOUT_TMP_0[12]\, RD11 => \DOUT_TMP_0[11]\, RD10 => 
        \DOUT_TMP_0[10]\, RD9 => \DOUT_TMP_0[9]\, RD8 => 
        \DOUT_TMP_0[8]\, RD7 => \DOUT_TMP_0[7]\, RD6 => 
        \DOUT_TMP_0[6]\, RD5 => \DOUT_TMP_0[5]\, RD4 => 
        \DOUT_TMP_0[4]\, RD3 => \DOUT_TMP_0[3]\, RD2 => 
        \DOUT_TMP_0[2]\, RD1 => \DOUT_TMP_0[1]\, RD0 => 
        \DOUT_TMP_0[0]\);
    
    rfd_tile_I_1_RNIB3001 : MX2
      port map(A => \DOUT_TMP[16]\, B => \DIN_REG1[16]\, S => 
        N_7_0, Y => hwdata_c(16));
    
    \rfd_tile_DIN_REG1[16]\ : DFN1
      port map(D => wdata(16), CLK => HCLK_c, Q => \DIN_REG1[16]\);
    
    \rfd_tile_WADDR_REG1[1]\ : DFN1
      port map(D => Waddr_vect_RNI0O455(1), CLK => HCLK_c, Q => 
        \WADDR_REG1[1]\);
    
    rfd_tile_I_1_RNIC3001 : MX2
      port map(A => \DOUT_TMP[17]\, B => \DIN_REG1[17]\, S => 
        N_7_0, Y => hwdata_c(17));
    
    \rfd_tile_RADDR_REG1_RNIQS1L_0[0]\ : NOR3C
      port map(A => I_5_1, B => I_5_0, C => I_5_5, Y => N_7);
    
    \rfd_tile_DIN_REG1[17]\ : DFN1
      port map(D => wdata(17), CLK => HCLK_c, Q => \DIN_REG1[17]\);
    
    \rfd_tile_0_DIN_REG1[4]\ : DFN1
      port map(D => wdata(22), CLK => HCLK_c, Q => \DIN_REG1[4]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    rfd_tile_I_1_RNI73001 : MX2
      port map(A => \DOUT_TMP_0[12]\, B => \DIN_REG1_0[12]\, S
         => N_7, Y => hwdata_c(12));
    
    \rfd_tile_DIN_REG1[7]\ : DFN1
      port map(D => wdata(7), CLK => HCLK_c, Q => \DIN_REG1_0[7]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity syncram_2pZ1 is

    port( hwdata_c            : out   std_logic_vector(31 downto 0);
          Raddr_vect_RNI4A0PH : in    std_logic_vector(0 to 0);
          Raddr_vect_RNICA1PH : in    std_logic_vector(1 to 1);
          Raddr_vect_RNIKA2PH : in    std_logic_vector(2 to 2);
          Raddr_vect_RNIE6Q5I : in    std_logic_vector(3 to 3);
          Raddr_vect_RNIIMQ5I : in    std_logic_vector(4 to 4);
          Waddr_vect_RNION355 : in    std_logic_vector(0 to 0);
          Waddr_vect_RNI0O455 : in    std_logic_vector(1 to 1);
          Waddr_vect_RNI394D5 : in    std_logic_vector(2 to 2);
          Waddr_vect_RNIJTNE5 : in    std_logic_vector(3 to 3);
          Waddr_vect_RNILLSP5 : in    std_logic_vector(4 to 4);
          wdata               : in    std_logic_vector(31 downto 0);
          HCLK_c              : in    std_logic;
          N_1_i_1             : in    std_logic;
          sEmpty_RNIE7T87     : in    std_logic;
          sEmpty_RNILSD08     : in    std_logic;
          sFull_RNIHL443      : in    std_logic;
          sFull_RNIU5GK1      : in    std_logic;
          syncram_2pZ1_GND    : in    std_logic;
          syncram_2pZ1_VCC    : in    std_logic;
          N_1_i_1_i           : in    std_logic
        );

end syncram_2pZ1;

architecture DEF_ARCH of syncram_2pZ1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component generic_syncram_2p_7_32_0
    port( wdata                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          Waddr_vect_RNILLSP5           : in    std_logic_vector(4 to 4) := (others => 'U');
          Waddr_vect_RNIJTNE5           : in    std_logic_vector(3 to 3) := (others => 'U');
          Waddr_vect_RNI394D5           : in    std_logic_vector(2 to 2) := (others => 'U');
          Waddr_vect_RNI0O455           : in    std_logic_vector(1 to 1) := (others => 'U');
          Waddr_vect_RNION355           : in    std_logic_vector(0 to 0) := (others => 'U');
          Raddr_vect_RNIIMQ5I           : in    std_logic_vector(4 to 4) := (others => 'U');
          Raddr_vect_RNIE6Q5I           : in    std_logic_vector(3 to 3) := (others => 'U');
          Raddr_vect_RNIKA2PH           : in    std_logic_vector(2 to 2) := (others => 'U');
          Raddr_vect_RNICA1PH           : in    std_logic_vector(1 to 1) := (others => 'U');
          Raddr_vect_RNI4A0PH           : in    std_logic_vector(0 to 0) := (others => 'U');
          hwdata_c                      : out   std_logic_vector(31 downto 0);
          N_1_i_1_i                     : in    std_logic := 'U';
          generic_syncram_2p_7_32_0_VCC : in    std_logic := 'U';
          generic_syncram_2p_7_32_0_GND : in    std_logic := 'U';
          sFull_RNIU5GK1                : in    std_logic := 'U';
          sFull_RNIHL443                : in    std_logic := 'U';
          sEmpty_RNILSD08               : in    std_logic := 'U';
          sEmpty_RNIE7T87               : in    std_logic := 'U';
          N_1_i_1                       : in    std_logic := 'U';
          HCLK_c                        : in    std_logic := 'U'
        );
  end component;

    signal \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : generic_syncram_2p_7_32_0
	Use entity work.generic_syncram_2p_7_32_0(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \inf.x0\ : generic_syncram_2p_7_32_0
      port map(wdata(31) => wdata(31), wdata(30) => wdata(30), 
        wdata(29) => wdata(29), wdata(28) => wdata(28), wdata(27)
         => wdata(27), wdata(26) => wdata(26), wdata(25) => 
        wdata(25), wdata(24) => wdata(24), wdata(23) => wdata(23), 
        wdata(22) => wdata(22), wdata(21) => wdata(21), wdata(20)
         => wdata(20), wdata(19) => wdata(19), wdata(18) => 
        wdata(18), wdata(17) => wdata(17), wdata(16) => wdata(16), 
        wdata(15) => wdata(15), wdata(14) => wdata(14), wdata(13)
         => wdata(13), wdata(12) => wdata(12), wdata(11) => 
        wdata(11), wdata(10) => wdata(10), wdata(9) => wdata(9), 
        wdata(8) => wdata(8), wdata(7) => wdata(7), wdata(6) => 
        wdata(6), wdata(5) => wdata(5), wdata(4) => wdata(4), 
        wdata(3) => wdata(3), wdata(2) => wdata(2), wdata(1) => 
        wdata(1), wdata(0) => wdata(0), Waddr_vect_RNILLSP5(4)
         => Waddr_vect_RNILLSP5(4), Waddr_vect_RNIJTNE5(3) => 
        Waddr_vect_RNIJTNE5(3), Waddr_vect_RNI394D5(2) => 
        Waddr_vect_RNI394D5(2), Waddr_vect_RNI0O455(1) => 
        Waddr_vect_RNI0O455(1), Waddr_vect_RNION355(0) => 
        Waddr_vect_RNION355(0), Raddr_vect_RNIIMQ5I(4) => 
        Raddr_vect_RNIIMQ5I(4), Raddr_vect_RNIE6Q5I(3) => 
        Raddr_vect_RNIE6Q5I(3), Raddr_vect_RNIKA2PH(2) => 
        Raddr_vect_RNIKA2PH(2), Raddr_vect_RNICA1PH(1) => 
        Raddr_vect_RNICA1PH(1), Raddr_vect_RNI4A0PH(0) => 
        Raddr_vect_RNI4A0PH(0), hwdata_c(31) => hwdata_c(31), 
        hwdata_c(30) => hwdata_c(30), hwdata_c(29) => 
        hwdata_c(29), hwdata_c(28) => hwdata_c(28), hwdata_c(27)
         => hwdata_c(27), hwdata_c(26) => hwdata_c(26), 
        hwdata_c(25) => hwdata_c(25), hwdata_c(24) => 
        hwdata_c(24), hwdata_c(23) => hwdata_c(23), hwdata_c(22)
         => hwdata_c(22), hwdata_c(21) => hwdata_c(21), 
        hwdata_c(20) => hwdata_c(20), hwdata_c(19) => 
        hwdata_c(19), hwdata_c(18) => hwdata_c(18), hwdata_c(17)
         => hwdata_c(17), hwdata_c(16) => hwdata_c(16), 
        hwdata_c(15) => hwdata_c(15), hwdata_c(14) => 
        hwdata_c(14), hwdata_c(13) => hwdata_c(13), hwdata_c(12)
         => hwdata_c(12), hwdata_c(11) => hwdata_c(11), 
        hwdata_c(10) => hwdata_c(10), hwdata_c(9) => hwdata_c(9), 
        hwdata_c(8) => hwdata_c(8), hwdata_c(7) => hwdata_c(7), 
        hwdata_c(6) => hwdata_c(6), hwdata_c(5) => hwdata_c(5), 
        hwdata_c(4) => hwdata_c(4), hwdata_c(3) => hwdata_c(3), 
        hwdata_c(2) => hwdata_c(2), hwdata_c(1) => hwdata_c(1), 
        hwdata_c(0) => hwdata_c(0), N_1_i_1_i => N_1_i_1_i, 
        generic_syncram_2p_7_32_0_VCC => syncram_2pZ1_VCC, 
        generic_syncram_2p_7_32_0_GND => syncram_2pZ1_GND, 
        sFull_RNIU5GK1 => sFull_RNIU5GK1, sFull_RNIHL443 => 
        sFull_RNIHL443, sEmpty_RNILSD08 => sEmpty_RNILSD08, 
        sEmpty_RNIE7T87 => sEmpty_RNIE7T87, N_1_i_1 => N_1_i_1, 
        HCLK_c => HCLK_c);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ2 is

    port( ready_i_0             : out   std_logic_vector(2 to 2);
          data_mem_wen_i_0      : out   std_logic_vector(2 to 2);
          data_ren              : in    std_logic_vector(2 to 2);
          Waddr_vect_RNI0O455   : out   std_logic_vector(1 to 1);
          Waddr_vect_RNILLSP5   : out   std_logic_vector(4 to 4);
          Waddr_vect_RNIJTNE5   : out   std_logic_vector(3 to 3);
          Waddr_vect_RNI394D5   : out   std_logic_vector(2 to 2);
          data_mem_ren_i_0_0    : in    std_logic;
          data_addr_r_0_iv_i_2  : in    std_logic_vector(5 to 5);
          data_addr_w_iv_i_4    : in    std_logic_vector(4 downto 0);
          Waddr_vect_RNION355   : out   std_logic_vector(0 to 0);
          data_wen              : in    std_logic_vector(2 to 2);
          data_addr_r_iv_i_a2_0 : in    std_logic_vector(4 to 4);
          data_addr_r_iv_i_a2_2 : out   std_logic_vector(4 to 4);
          HRESETn_c             : in    std_logic;
          HCLK_c                : in    std_logic;
          N_67                  : out   std_logic;
          N_166                 : in    std_logic;
          N_75                  : out   std_logic;
          N_59                  : out   std_logic;
          N_51                  : out   std_logic;
          N_43                  : out   std_logic;
          N_152                 : in    std_logic;
          N_128                 : in    std_logic;
          N_136                 : in    std_logic;
          N_144                 : in    std_logic;
          sEmpty_RNIE7T87       : out   std_logic;
          N_160                 : in    std_logic;
          N_77                  : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ2;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ2 is 

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_12, \data_mem_addr_w_2[1]\, \data_mem_addr_w_2[0]\, 
        N_4, \data_mem_addr_w_2[3]\, \DWACT_FINC_E[0]\, N_12_0, 
        \data_mem_addr_r_2[1]\, \data_mem_addr_r_2[0]\, N_4_0, 
        \data_mem_addr_r_2[3]\, \DWACT_FINC_E_0[0]\, 
        \data_mem_ren_i_0[2]\, un7_sempty_s_4, un7_sempty_s_1, 
        un7_sempty_s_0, un7_sempty_s_2, \sEmpty_RNO_6\, 
        \sEmpty_RNO_7\, \un10_raddr_vect_s[1]\, \sEmpty_RNO_5\, 
        \un10_raddr_vect_s[0]\, un5_sfull_s_4_2, 
        \un8_waddr_vect_s[3]\, sFull_RNO_8_0, un5_sfull_s_4_1, 
        \un8_waddr_vect_s[1]\, sFull_RNO_5_2, un5_sfull_s_4_0, 
        \un8_waddr_vect_s[0]\, ADD_7x7_fast_I23_Y_0_o2_0, N165_1, 
        N_89_i, N_109, ADD_5x5_fast_I11_Y_i_a2_1, 
        ADD_5x5_fast_I11_Y_i_a2_0, N_17, \data_mem_addr_r_2[2]\, 
        \data_mem_addr_w_2[2]\, SUM2_0_0, ADD_5x5_fast_I11_Y_0, 
        N80, un1_waddr_vect_slto3_0, un2_raddr_vect_slto3_0, 
        N_159, N_143, N_135, N_127, N_151, \un117_ready1[4]\, 
        N_87, CO1_tz, N_12_1, N_18, I11_un1_Y, N81, N77, N98, 
        un5_sfull_s_4, Waddr_vect_n4, \data_mem_addr_w_2[4]\, 
        Waddr_vect_14_0, N_58_i_0, Waddr_vect_c2, Waddr_vect_n3, 
        sFull_RNO_9, \sFull\, ADD_7x7_fast_I19_Y_i_a2_0_206, 
        N_9_i, N_105_1, Waddr_vect_n2, Waddr_vect_c1_i_0, 
        \sEmpty\, un1_sempty_s, sEmpty_RNO_10, un2_raddr_vect_s, 
        I_5_16, \un10_raddr_vect_s[2]\, I_9_16, 
        \un10_raddr_vect_s[3]\, I_13_16, \un10_raddr_vect_s[4]\, 
        I_20_8, I_5_15, I_13_15, \data_mem_addr_r_2[4]\, 
        \data_mem_wen_i_0[2]\, Waddr_vect_e1, Waddr_vect_n1_i, 
        Waddr_vect_e4, I_20_7, I_9_15, Waddr_vect_e3, 
        Waddr_vect_e0, N_85_i, N_24, N_75_0, \un132_ready1[4]\, 
        I8_un1_Y, \un132_ready0_1[4]\, \un117_ready0[4]\, N_6, 
        \un132_ready0[4]\, un119_readylto4, un134_ready, 
        un126_ready, N_198, N107, N161, N_197, \un132_ready1[5]\, 
        N_16_i_i_0, N_196, N_13, un2_raddr_vect_slto1, 
        Waddr_vect_e2, N_9, N_13_0, N_12_2, N_11, N_8, N_10, 
        N_9_0, N_7, N_4_1, N_5, N_6_0, N_9_1, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 

    data_mem_wen_i_0(2) <= \data_mem_wen_i_0[2]\;

    un117_ready_1_1_0_CO1_tz : AO18
      port map(A => N_105_1, B => \data_mem_addr_w_2[2]\, C => 
        \data_mem_addr_r_2[2]\, Y => CO1_tz);
    
    sFull : DFN1C0
      port map(D => sFull_RNO_9, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => \sFull\);
    
    un117_ready_1_1_0_SUM2_0 : AX1C
      port map(A => N_87, B => CO1_tz, C => SUM2_0_0, Y => 
        \un117_ready1[4]\);
    
    \ready_gen.un126_ready_0_I_11\ : OA1
      port map(A => N_13_0, B => N_12_2, C => N_11, Y => 
        un126_ready);
    
    \Waddr_vect_RNO[0]\ : AXOI5
      port map(A => N_58_i_0, B => \data_mem_wen_i_0[2]\, C => 
        \data_mem_addr_w_2[0]\, Y => Waddr_vect_e0);
    
    sFull_RNO_8 : AX1E
      port map(A => N_58_i_0, B => I_20_7, C => 
        \data_mem_addr_r_2[4]\, Y => sFull_RNO_8_0);
    
    un117_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0_0 : AO1C
      port map(A => \data_mem_addr_r_2[2]\, B => 
        \data_mem_addr_w_2[2]\, C => N_109, Y => 
        ADD_5x5_fast_I11_Y_i_a2_0);
    
    sFull_RNO_6 : OR2A
      port map(A => N_58_i_0, B => \data_mem_addr_w_2[0]\, Y => 
        \un8_waddr_vect_s[0]\);
    
    \Raddr_vect_RNIVJ63[1]\ : OR2B
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \data_mem_addr_r_2[0]\, Y => un2_raddr_vect_slto1);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_2[0]\);
    
    \Raddr_vect_RNI53FB1[0]\ : MX2
      port map(A => \un117_ready1[4]\, B => \un117_ready0[4]\, S
         => \data_mem_addr_r_2[0]\, Y => un119_readylto4);
    
    un132_ready_1_16_ADD_5x5_fast_I11_Y_0 : AO1
      port map(A => N80, B => N_109, C => N_89_i, Y => 
        ADD_5x5_fast_I11_Y_0);
    
    un132_ready_0_0_0_ADD_7x7_fast_I23_Y_0_o2_0 : AO1A
      port map(A => N165_1, B => N_89_i, C => N_109, Y => 
        ADD_7x7_fast_I23_Y_0_o2_0);
    
    \Waddr_vect_RNO[3]\ : MX2B
      port map(A => \data_mem_addr_w_2[3]\, B => Waddr_vect_n3, S
         => \data_mem_wen_i_0[2]\, Y => Waddr_vect_e3);
    
    \Waddr_vect_RNI394D5[2]\ : NOR3C
      port map(A => data_addr_w_iv_i_4(2), B => N_143, C => N_144, 
        Y => Waddr_vect_RNI394D5(2));
    
    \Raddr_vect_RNI8ULN5[0]\ : AOI1
      port map(A => N_197, B => N_196, C => N_198, Y => 
        un134_ready);
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \data_mem_addr_r_2[0]\, Y => N_12_0);
    
    \Waddr_vect_RNION355[0]\ : NOR3C
      port map(A => data_addr_w_iv_i_4(0), B => N_159, C => N_160, 
        Y => Waddr_vect_RNION355(0));
    
    \Waddr_vect_RNIPN791[0]\ : OR3A
      port map(A => \data_mem_wen_i_0[2]\, B => N_166, C => 
        \data_mem_addr_w_2[0]\, Y => N_159);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_w_2[0]\, B => 
        \data_mem_addr_w_2[1]\, Y => I_5_15);
    
    un132_ready_1_16_ADD_5x5_fast_I8_un1_Y : NOR2B
      port map(A => N81, B => N77, Y => I8_un1_Y);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => un7_sempty_s_1, B => un7_sempty_s_0, C => 
        un7_sempty_s_2, Y => un7_sempty_s_4);
    
    un132_ready_0_0_0_ADD_7x7_fast_I33_Y_0_i_x2 : AX1E
      port map(A => N_24, B => ADD_7x7_fast_I23_Y_0_o2_0, C => 
        N_75_0, Y => N_16_i_i_0);
    
    \Raddr_vect_RNI5KRC[4]\ : NOR2B
      port map(A => I_9_16, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[2]\);
    
    \Waddr_vect_RNIT7891[4]\ : OR3A
      port map(A => \data_mem_wen_i_0[2]\, B => N_166, C => 
        \data_mem_addr_w_2[4]\, Y => N_127);
    
    un117_ready_0_0_0_ADD_5x5_fast_I18_Y_0 : XNOR2
      port map(A => N_6, B => N_89_i, Y => \un117_ready0[4]\);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_r_2[0]\, B => 
        \data_mem_addr_r_2[1]\, C => \data_mem_addr_r_2[2]\, Y
         => N_9);
    
    un117_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3 : NOR2
      port map(A => N_9_i, B => \data_mem_addr_r_2[2]\, Y => N_17);
    
    \Raddr_vect_RNI7073[2]\ : XNOR2
      port map(A => \data_mem_addr_w_2[2]\, B => 
        \data_mem_addr_r_2[2]\, Y => N_85_i);
    
    \ready_gen.un126_ready_0_I_4\ : OR2A
      port map(A => \data_mem_addr_r_2[4]\, B => 
        \data_mem_addr_w_2[4]\, Y => N_7);
    
    \Waddr_vect_RNO[4]\ : MX2B
      port map(A => \data_mem_addr_w_2[4]\, B => Waddr_vect_n4, S
         => \data_mem_wen_i_0[2]\, Y => Waddr_vect_e4);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_2[1]\);
    
    sFull_RNO_7 : OR2B
      port map(A => I_13_15, B => N_58_i_0, Y => 
        \un8_waddr_vect_s[3]\);
    
    \Raddr_vect_RNIB3352[1]\ : OR2
      port map(A => \data_mem_ren_i_0[2]\, B => 
        \data_mem_addr_r_2[1]\, Y => N_67);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_9_1, B => \data_mem_addr_w_2[3]\, Y => 
        I_13_15);
    
    GND_i : GND
      port map(Y => \GND\);
    
    sEmpty_RNO_7 : XNOR2
      port map(A => \un10_raddr_vect_s[4]\, B => 
        \data_mem_addr_w_2[4]\, Y => \sEmpty_RNO_7\);
    
    un117_ready_0_0_0_ADD_5x5_fast_I11_Y_i : OR2B
      port map(A => N_13, B => N_12_1, Y => N_6);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Raddr_vect_RNI5O63[1]\ : NOR2A
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \data_mem_addr_w_2[1]\, Y => N_105_1);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_w_2[0]\, B => 
        \data_mem_addr_w_2[1]\, C => \data_mem_addr_w_2[2]\, Y
         => N_9_1);
    
    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \data_mem_addr_w_2[1]\, B => 
        \data_mem_addr_w_2[0]\, C => N_58_i_0, Y => 
        Waddr_vect_n1_i);
    
    un117_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_1 : OR2
      port map(A => ADD_5x5_fast_I11_Y_i_a2_0, B => N_17, Y => 
        ADD_5x5_fast_I11_Y_i_a2_1);
    
    \Raddr_vect[2]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[2]\, Q => 
        \data_mem_addr_r_2[2]\);
    
    un117_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2 : OR2
      port map(A => ADD_5x5_fast_I11_Y_i_a2_1, B => N_18, Y => 
        N_12_1);
    
    un132_ready_1_16_ADD_5x5_fast_I1_G0N : AO1C
      port map(A => \data_mem_addr_w_2[2]\, B => 
        \data_mem_addr_r_2[2]\, C => N_87, Y => N80);
    
    \Waddr_vect_RNIS3891[3]\ : OR3A
      port map(A => \data_mem_wen_i_0[2]\, B => N_166, C => 
        \data_mem_addr_w_2[3]\, Y => N_135);
    
    \Raddr_vect_RNIGJ408[0]\ : MX2
      port map(A => un119_readylto4, B => un134_ready, S => 
        un126_ready, Y => ready_i_0(2));
    
    \Raddr_vect_RNI9873_0[3]\ : OR2A
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \data_mem_addr_r_2[3]\, Y => N_109);
    
    \Waddr_vect_RNO_0[4]\ : XAI1A
      port map(A => \data_mem_addr_w_2[4]\, B => Waddr_vect_14_0, 
        C => N_58_i_0, Y => Waddr_vect_n4);
    
    un132_ready_1_16_ADD_5x5_fast_I0_CO1 : NOR2
      port map(A => N_105_1, B => N_85_i, Y => N77);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    sEmpty_RNIT8VB4 : NOR3C
      port map(A => N_77, B => data_addr_r_iv_i_a2_0(4), C => 
        \data_mem_ren_i_0[2]\, Y => data_addr_r_iv_i_a2_2(4));
    
    sEmpty_RNO : AO1A
      port map(A => data_ren(2), B => un7_sempty_s_4, C => 
        un1_sempty_s, Y => sEmpty_RNO_10);
    
    \Waddr_vect[3]\ : DFN1C0
      port map(D => Waddr_vect_e3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_2[3]\);
    
    \Raddr_vect_RNIAV252[0]\ : OR2
      port map(A => \data_mem_ren_i_0[2]\, B => 
        \data_mem_addr_r_2[0]\, Y => N_75);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_w_2[1]\, B => 
        \data_mem_addr_w_2[0]\, Y => N_12);
    
    sEmpty_RNO_3 : XA1A
      port map(A => \data_mem_addr_w_2[0]\, B => 
        \un10_raddr_vect_s[0]\, C => data_wen(2), Y => 
        un7_sempty_s_0);
    
    \Waddr_vect_RNIUG18[4]\ : AO1B
      port map(A => un1_waddr_vect_slto3_0, B => 
        Waddr_vect_c1_i_0, C => \data_mem_addr_w_2[4]\, Y => 
        N_58_i_0);
    
    un6_waddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \DWACT_FINC_E[0]\, Y => N_4);
    
    \Raddr_vect_RNI5G18[4]\ : AO1B
      port map(A => un2_raddr_vect_slto3_0, B => 
        un2_raddr_vect_slto1, C => \data_mem_addr_r_2[4]\, Y => 
        un2_raddr_vect_s);
    
    \Waddr_vect[4]\ : DFN1C0
      port map(D => Waddr_vect_e4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_2[4]\);
    
    sFull_RNO : OA1
      port map(A => \sFull\, B => un5_sfull_s_4, C => data_ren(2), 
        Y => sFull_RNO_9);
    
    \Raddr_vect_RNIA03G[4]\ : NOR2B
      port map(A => I_20_8, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[4]\);
    
    \ready_gen.un126_ready_0_I_9\ : AO1C
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \data_mem_addr_r_2[3]\, C => N_7, Y => N_12_2);
    
    sFull_RNO_2 : XA1B
      port map(A => \data_mem_addr_r_2[0]\, B => 
        \un8_waddr_vect_s[0]\, C => data_wen(2), Y => 
        un5_sfull_s_4_0);
    
    \ready_gen.un126_ready_0_I_7\ : AO1C
      port map(A => \data_mem_addr_w_2[2]\, B => 
        \data_mem_addr_r_2[2]\, C => N_4_1, Y => N_10);
    
    un132_ready_0_0_0_ADD_7x7_fast_I32_Y_0 : AX1A
      port map(A => N165_1, B => N80, C => \un132_ready0_1[4]\, Y
         => \un132_ready0[4]\);
    
    \Waddr_vect_RNO_0[2]\ : XAI1A
      port map(A => \data_mem_addr_w_2[2]\, B => 
        Waddr_vect_c1_i_0, C => N_58_i_0, Y => Waddr_vect_n2);
    
    \ready_gen.un126_ready_0_I_5\ : AO1C
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \data_mem_addr_w_2[1]\, C => N_6_0, Y => N_8);
    
    \ready_gen.un126_ready_0_I_3\ : NOR2A
      port map(A => \data_mem_addr_r_2[0]\, B => 
        \data_mem_addr_w_2[0]\, Y => N_6_0);
    
    un132_ready_1_16_ADD_5x5_fast_I16_Y_0 : AX1E
      port map(A => I11_un1_Y, B => ADD_5x5_fast_I11_Y_0, C => 
        N_75_0, Y => \un132_ready1[5]\);
    
    \Raddr_vect[0]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[2]\, Q => 
        \data_mem_addr_r_2[0]\);
    
    sFull_RNIDVR9 : NOR2
      port map(A => \sFull\, B => data_wen(2), Y => 
        \data_mem_wen_i_0[2]\);
    
    \Waddr_vect_RNO_0[3]\ : XAI1
      port map(A => \data_mem_addr_w_2[3]\, B => Waddr_vect_c2, C
         => N_58_i_0, Y => Waddr_vect_n3);
    
    \ready_gen.un126_ready_0_I_6\ : OA1A
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \data_mem_addr_r_2[3]\, C => N_5, Y => N_9_0);
    
    \Waddr_vect_RNI0O455[1]\ : NOR3C
      port map(A => data_addr_w_iv_i_4(1), B => N_151, C => N_152, 
        Y => Waddr_vect_RNI0O455(1));
    
    un132_ready_1_16_ADD_5x5_fast_I1_P0N : OR3A
      port map(A => \data_mem_addr_r_2[2]\, B => 
        \data_mem_addr_w_2[2]\, C => N_87, Y => N81);
    
    sEmpty_RNIBNF32 : OR2
      port map(A => \sEmpty\, B => data_ren(2), Y => 
        \data_mem_ren_i_0[2]\);
    
    \Raddr_vect_RNI4OK9[0]\ : NOR2A
      port map(A => un2_raddr_vect_s, B => \data_mem_addr_r_2[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_12_0, B => \data_mem_addr_r_2[2]\, Y => 
        I_9_16);
    
    \sEmpty_RNIE7T87\ : NOR3B
      port map(A => \data_mem_ren_i_0[2]\, B => 
        data_addr_r_0_iv_i_2(5), C => data_mem_ren_i_0_0, Y => 
        sEmpty_RNIE7T87);
    
    \Raddr_vect_RNIBG73[4]\ : XNOR2
      port map(A => \data_mem_addr_w_2[4]\, B => 
        \data_mem_addr_r_2[4]\, Y => N_89_i);
    
    \Waddr_vect_RNIRV791[2]\ : OR3A
      port map(A => \data_mem_wen_i_0[2]\, B => N_166, C => 
        \data_mem_addr_w_2[2]\, Y => N_143);
    
    \Waddr_vect_RNIQR791[1]\ : OR3A
      port map(A => \data_mem_wen_i_0[2]\, B => N_166, C => 
        \data_mem_addr_w_2[1]\, Y => N_151);
    
    sFull_RNO_3 : XA1
      port map(A => \data_mem_addr_r_2[3]\, B => 
        \un8_waddr_vect_s[3]\, C => sFull_RNO_8_0, Y => 
        un5_sfull_s_4_2);
    
    un8_raddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_r_2[0]\, B => 
        \data_mem_addr_r_2[1]\, C => \data_mem_addr_r_2[2]\, Y
         => \DWACT_FINC_E_0[0]\);
    
    \ready_gen.un126_ready_0_I_1\ : OR2A
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \data_mem_addr_w_2[1]\, Y => N_4_1);
    
    \Waddr_vect_RNO_1[4]\ : OR2B
      port map(A => Waddr_vect_c2, B => \data_mem_addr_w_2[3]\, Y
         => Waddr_vect_14_0);
    
    \Raddr_vect_RNIC7352[2]\ : OR2
      port map(A => \data_mem_ren_i_0[2]\, B => 
        \data_mem_addr_r_2[2]\, Y => N_59);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Raddr_vect_RNI9873[3]\ : XNOR2
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \data_mem_addr_r_2[3]\, Y => N_87);
    
    \Raddr_vect_RNI3473[3]\ : NOR2
      port map(A => \data_mem_addr_r_2[3]\, B => 
        \data_mem_addr_r_2[2]\, Y => un2_raddr_vect_slto3_0);
    
    un132_ready_0_0_0_ADD_7x7_fast_I23_Y_0 : OR2A
      port map(A => N_75_0, B => \un117_ready0[4]\, Y => N161);
    
    un6_waddr_vect_s_I_20 : XOR2
      port map(A => N_4, B => \data_mem_addr_w_2[4]\, Y => I_20_7);
    
    \Raddr_vect[1]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[2]\, Q => 
        \data_mem_addr_r_2[1]\);
    
    un132_ready_0_0_0_ADD_7x7_fast_I19_Y_i_a2_0_206 : NOR2A
      port map(A => \data_mem_addr_w_2[2]\, B => 
        \data_mem_addr_r_2[2]\, Y => 
        ADD_7x7_fast_I19_Y_i_a2_0_206);
    
    sEmpty_RNO_6 : XNOR2
      port map(A => \un10_raddr_vect_s[3]\, B => 
        \data_mem_addr_w_2[3]\, Y => \sEmpty_RNO_6\);
    
    \Raddr_vect_RNIBG73_0[4]\ : NOR2A
      port map(A => \data_mem_addr_r_2[4]\, B => 
        \data_mem_addr_w_2[4]\, Y => N_75_0);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_9, B => \data_mem_addr_r_2[3]\, Y => 
        I_13_16);
    
    \ready_gen.un126_ready_0_I_8\ : OR2A
      port map(A => \data_mem_addr_w_2[4]\, B => 
        \data_mem_addr_r_2[4]\, Y => N_11);
    
    \Waddr_vect_RNO[2]\ : MX2B
      port map(A => \data_mem_addr_w_2[2]\, B => Waddr_vect_n2, S
         => \data_mem_wen_i_0[2]\, Y => Waddr_vect_e2);
    
    sFull_RNO_0 : NOR3C
      port map(A => un5_sfull_s_4_1, B => un5_sfull_s_4_0, C => 
        un5_sfull_s_4_2, Y => un5_sfull_s_4);
    
    sEmpty_RNO_2 : XA1A
      port map(A => \data_mem_addr_w_2[1]\, B => 
        \un10_raddr_vect_s[1]\, C => \sEmpty_RNO_5\, Y => 
        un7_sempty_s_1);
    
    \Raddr_vect_RNISJHJ1[0]\ : MX2C
      port map(A => \un132_ready1[4]\, B => \un132_ready0[4]\, S
         => \data_mem_addr_r_2[0]\, Y => N_196);
    
    sEmpty_RNO_4 : NOR2B
      port map(A => \sEmpty_RNO_6\, B => \sEmpty_RNO_7\, Y => 
        un7_sempty_s_2);
    
    sFull_RNO_5 : AX1E
      port map(A => N_58_i_0, B => I_9_15, C => 
        \data_mem_addr_r_2[2]\, Y => sFull_RNO_5_2);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_r_2[0]\, B => 
        \data_mem_addr_r_2[1]\, Y => I_5_16);
    
    \Waddr_vect_RNIJTNE5[3]\ : NOR3C
      port map(A => data_addr_w_iv_i_4(3), B => N_135, C => N_136, 
        Y => Waddr_vect_RNIJTNE5(3));
    
    un117_ready_1_1_0_SUM2_0_0 : XNOR2
      port map(A => N_109, B => N_89_i, Y => SUM2_0_0);
    
    \Waddr_vect_RNI9K63[0]\ : OR2B
      port map(A => \data_mem_addr_w_2[1]\, B => 
        \data_mem_addr_w_2[0]\, Y => Waddr_vect_c1_i_0);
    
    un132_ready_1_16_ADD_5x5_fast_I15_Y_0 : AX1A
      port map(A => I8_un1_Y, B => N80, C => \un132_ready0_1[4]\, 
        Y => \un132_ready1[4]\);
    
    \ready_gen.un126_ready_0_I_10\ : OA1A
      port map(A => N_8, B => N_10, C => N_9_0, Y => N_13_0);
    
    sEmpty : DFN1P0
      port map(D => sEmpty_RNO_10, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \sEmpty\);
    
    \Waddr_vect_RNO[1]\ : MX2B
      port map(A => \data_mem_addr_w_2[1]\, B => Waddr_vect_n1_i, 
        S => \data_mem_wen_i_0[2]\, Y => Waddr_vect_e1);
    
    \Raddr_vect_RNI448B[4]\ : NOR2B
      port map(A => I_5_16, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[1]\);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_2[2]\);
    
    un132_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1 : OA1B
      port map(A => ADD_7x7_fast_I19_Y_i_a2_0_206, B => N_87, C
         => N_9_i, Y => N165_1);
    
    un6_waddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_w_2[0]\, B => 
        \data_mem_addr_w_2[1]\, C => \data_mem_addr_w_2[2]\, Y
         => \DWACT_FINC_E[0]\);
    
    un117_ready_0_0_0_ADD_5x5_fast_I9_Y_i_o2 : AO18
      port map(A => \data_mem_addr_w_2[1]\, B => 
        \data_mem_addr_r_2[1]\, C => \data_mem_addr_w_2[0]\, Y
         => N_9_i);
    
    un132_ready_0_0_0_ADD_7x7_fast_I23_Y_0_a4_0 : AO1A
      port map(A => N165_1, B => N80, C => N_89_i, Y => N_24);
    
    sFull_RNO_1 : XA1
      port map(A => \data_mem_addr_r_2[1]\, B => 
        \un8_waddr_vect_s[1]\, C => sFull_RNO_5_2, Y => 
        un5_sfull_s_4_1);
    
    \Waddr_vect_RNILLSP5[4]\ : NOR3C
      port map(A => data_addr_w_iv_i_4(4), B => N_127, C => N_128, 
        Y => Waddr_vect_RNILLSP5(4));
    
    un132_ready_1_16_ADD_5x5_fast_I10_Y : OR2B
      port map(A => I11_un1_Y, B => N_75_0, Y => N107);
    
    un132_ready_0_0_0_ADD_7x7_fast_I32_Y_0_1 : XOR2
      port map(A => N_109, B => N_89_i, Y => \un132_ready0_1[4]\);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[2]\, Q => 
        \data_mem_addr_r_2[3]\);
    
    sFull_RNO_4 : OR2B
      port map(A => I_5_15, B => N_58_i_0, Y => 
        \un8_waddr_vect_s[1]\);
    
    \Raddr_vect_RNI78FE[4]\ : NOR2B
      port map(A => I_13_16, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    sEmpty_RNO_5 : XNOR2
      port map(A => \un10_raddr_vect_s[2]\, B => 
        \data_mem_addr_w_2[2]\, Y => \sEmpty_RNO_5\);
    
    \Waddr_vect_RNID473[3]\ : NOR2
      port map(A => \data_mem_addr_w_2[3]\, B => 
        \data_mem_addr_w_2[2]\, Y => un1_waddr_vect_slto3_0);
    
    un117_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3_0 : NOR2A
      port map(A => \data_mem_addr_w_2[2]\, B => N_9_i, Y => N_18);
    
    un132_ready_1_16_ADD_5x5_fast_I11_un1_Y : OR3C
      port map(A => N81, B => N77, C => N98, Y => I11_un1_Y);
    
    \ready_gen.un126_ready_0_I_2\ : OR2A
      port map(A => \data_mem_addr_w_2[2]\, B => 
        \data_mem_addr_r_2[2]\, Y => N_5);
    
    \Raddr_vect_RNI245L1[0]\ : MX2C
      port map(A => N107, B => N161, S => \data_mem_addr_r_2[0]\, 
        Y => N_198);
    
    un8_raddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_r_2[3]\, B => 
        \DWACT_FINC_E_0[0]\, Y => N_4_0);
    
    \Waddr_vect_RNIF4Q4[2]\ : NOR2A
      port map(A => \data_mem_addr_w_2[2]\, B => 
        Waddr_vect_c1_i_0, Y => Waddr_vect_c2);
    
    \Raddr_vect_RNIA6VE2[0]\ : MX2C
      port map(A => \un132_ready1[5]\, B => N_16_i_i_0, S => 
        \data_mem_addr_r_2[0]\, Y => N_197);
    
    \Raddr_vect[4]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[2]\, Q => 
        \data_mem_addr_r_2[4]\);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_12, B => \data_mem_addr_w_2[2]\, Y => 
        I_9_15);
    
    un117_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0 : OR2A
      port map(A => \data_mem_addr_r_2[3]\, B => 
        \data_mem_addr_w_2[3]\, Y => N_13);
    
    sEmpty_RNO_1 : NOR2B
      port map(A => \sEmpty\, B => data_wen(2), Y => un1_sempty_s);
    
    \Raddr_vect_RNIDB352[3]\ : OR2
      port map(A => \data_mem_ren_i_0[2]\, B => 
        \data_mem_addr_r_2[3]\, Y => N_51);
    
    \Raddr_vect_RNIEF352[4]\ : OR2
      port map(A => \data_mem_ren_i_0[2]\, B => 
        \data_mem_addr_r_2[4]\, Y => N_43);
    
    un132_ready_1_16_ADD_5x5_fast_I2_P0N : OR2B
      port map(A => N_109, B => N_89_i, Y => N98);
    
    un8_raddr_vect_s_I_20 : XOR2
      port map(A => N_4_0, B => \data_mem_addr_r_2[4]\, Y => 
        I_20_8);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ5 is

    port( time_mem_wen_i_0_0 : in    std_logic;
          Waddr_vect_RNINV58 : out   std_logic_vector(2 to 2);
          Waddr_vect_RNILN58 : out   std_logic_vector(0 to 0);
          Raddr_vect_RNI8J9L : out   std_logic_vector(2 to 2);
          time_mem_ren_i_0   : out   std_logic_vector(1 to 1);
          time_wen           : in    std_logic_vector(1 to 1);
          time_ren           : in    std_logic_vector(1 to 1);
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic;
          N_146              : out   std_logic;
          N_162              : out   std_logic;
          N_113              : out   std_logic;
          N_122              : out   std_logic;
          sFull_RNIPQBB_0    : out   std_logic;
          N_62               : out   std_logic;
          N_70               : out   std_logic;
          sEmpty_RNI5EFO_0   : out   std_logic;
          N_33               : out   std_logic;
          N_29               : out   std_logic
        );

end lpp_waveform_fifo_ctrlZ5;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ5 is 

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \time_mem_addr_r_1[5]\, \Raddr_vect[2]_net_1\, 
        \Raddr_vect[3]_net_1\, \DWACT_FINC_E[0]\, 
        \time_mem_addr_w_1[5]\, \Waddr_vect[2]_net_1\, 
        \Waddr_vect[3]_net_1\, \DWACT_FINC_E_0[0]\, N_7, 
        \time_mem_addr_r_1[1]\, \time_mem_addr_r_1[0]\, N_7_0, 
        \time_mem_addr_w_1[1]\, \time_mem_addr_w_1[0]\, 
        un5_sfull_s_2, \un8_waddr_vect_s[3]\, un5_sfull_s_1, 
        \un8_waddr_vect_s[1]\, sFull_RNO_5_0, un5_sfull_s_0, 
        \un8_waddr_vect_s[0]\, un7_sempty_s_3, sEmpty_RNO_3_1, 
        sEmpty_RNO_4_1, un7_sempty_s_0, un7_sempty_s_2, 
        \un10_raddr_vect_s[3]\, \un10_raddr_vect_s[0]\, 
        un1_waddr_vect_slt3, un5_sfull_s, un2_raddr_vect_slt3, 
        Raddr_vect_n3, Raddr_vect_7_0, Waddr_vect_n3, 
        Waddr_vect_15_0, Raddr_vect_n2, un2_raddr_vect_s, 
        Raddr_vect_n2_tz, Waddr_vect_n2, un1_waddr_vect_s, 
        Waddr_vect_n2_tz, \time_mem_ren_i_0[1]\, 
        \time_mem_addr_r_1[3]\, N_167, I_9_10, Raddr_vect_n1_i, 
        Raddr_vect_e2, Raddr_vect_e1, Raddr_vect_e0, I_13_10, 
        I_9_9, I_5_10, Waddr_vect_n1_i, Waddr_vect_e2, 
        \time_mem_wen_i_0[1]\, Waddr_vect_e1, Waddr_vect_e0, 
        I_13_9, I_5_9, \sFull_RNO_2\, \sFull\, \sEmpty_RNO_2\, 
        un2_sempty_s, \sEmpty\, \time_mem_addr_w_1[3]\, N_4, 
        N_4_0, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    time_mem_ren_i_0(1) <= \time_mem_ren_i_0[1]\;

    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_w_1[1]\, B => 
        \time_mem_addr_w_1[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_w_1[0]\, B => 
        \time_mem_addr_w_1[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        N_4);
    
    sFull_RNIPQBB_1 : NOR2
      port map(A => \time_mem_addr_w_1[5]\, B => N_167, Y => 
        N_122);
    
    \Raddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_r_1[1]\, B => 
        \time_mem_addr_r_1[0]\, C => un2_raddr_vect_s, Y => 
        Raddr_vect_n1_i);
    
    sEmpty_RNI5EFO_1 : NOR2
      port map(A => \time_mem_ren_i_0[1]\, B => 
        \time_mem_addr_r_1[5]\, Y => N_33);
    
    un36_mem_addr_wen_I_8 : OR2B
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_1[5]\);
    
    un36_mem_addr_wen_I_16 : NOR2B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \Waddr_vect[2]_net_1\, Y => \DWACT_FINC_E_0[0]\);
    
    \Waddr_vect_RNI0PG9[1]\ : OR3
      port map(A => \time_mem_addr_w_1[0]\, B => 
        \time_mem_addr_w_1[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        un1_waddr_vect_slt3);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_w_1[1]\, B => 
        \time_mem_addr_w_1[0]\, Y => N_7_0);
    
    sEmpty_RNO : AO1
      port map(A => un7_sempty_s_3, B => un7_sempty_s_2, C => 
        un2_sempty_s, Y => \sEmpty_RNO_2\);
    
    \Raddr_vect[1]\ : DFN1C0
      port map(D => Raddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_1[1]\);
    
    \Waddr_vect[3]\ : DFN1E0C0
      port map(D => Waddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_wen_i_0[1]\, Q => 
        \Waddr_vect[3]_net_1\);
    
    sEmpty_RNI5EFO : OR2A
      port map(A => \DWACT_FINC_E[0]\, B => \time_mem_ren_i_0[1]\, 
        Y => N_29);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_7, B => \Raddr_vect[2]_net_1\, Y => I_9_10);
    
    \Raddr_vect_RNI7F9L[1]\ : OR2
      port map(A => \time_mem_ren_i_0[1]\, B => 
        \time_mem_addr_r_1[1]\, Y => N_62);
    
    sEmpty : DFN1P0
      port map(D => \sEmpty_RNO_2\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \sEmpty\);
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => \time_mem_wen_i_0[1]\, 
        C => \time_mem_addr_w_1[0]\, Y => Waddr_vect_e0);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Waddr_vect[2]_net_1\);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \time_mem_addr_w_1[1]\, 
        S => \time_mem_wen_i_0[1]\, Y => Waddr_vect_e1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Waddr_vect_RNO_0[2]\ : OR2B
      port map(A => un1_waddr_vect_s, B => Waddr_vect_n2_tz, Y
         => Waddr_vect_n2);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_w_1[0]\, B => 
        \time_mem_addr_w_1[1]\, Y => I_5_9);
    
    \Raddr_vect_RNO_0[2]\ : OR2B
      port map(A => un2_raddr_vect_s, B => Raddr_vect_n2_tz, Y
         => Raddr_vect_n2);
    
    sFull_RNIM805_0 : OR2A
      port map(A => time_mem_wen_i_0_0, B => 
        \time_mem_wen_i_0[1]\, Y => N_167);
    
    sFull_RNIPQBB : OR2A
      port map(A => \DWACT_FINC_E_0[0]\, B => N_167, Y => N_113);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => Raddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_ren_i_0[1]\, Q => 
        \Raddr_vect[3]_net_1\);
    
    \sFull_RNIPQBB_0\ : OR2
      port map(A => \time_mem_addr_w_1[3]\, B => N_167, Y => 
        sFull_RNIPQBB_0);
    
    sEmpty_RNO_2 : NOR2B
      port map(A => time_wen(1), B => \sEmpty\, Y => un2_sempty_s);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_4, B => \Waddr_vect[3]_net_1\, Y => I_13_9);
    
    un31_mem_addr_ren_I_5 : XOR2
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_1[3]\);
    
    sFull_RNO : AO1
      port map(A => time_ren(1), B => \sFull\, C => un5_sfull_s, 
        Y => \sFull_RNO_2\);
    
    \Raddr_vect_RNO[0]\ : AXOI7
      port map(A => un2_raddr_vect_s, B => \time_mem_ren_i_0[1]\, 
        C => \time_mem_addr_r_1[0]\, Y => Raddr_vect_e0);
    
    \Raddr_vect_RNO[1]\ : MX2A
      port map(A => Raddr_vect_n1_i, B => \time_mem_addr_r_1[1]\, 
        S => \time_mem_ren_i_0[1]\, Y => Raddr_vect_e1);
    
    sFull_RNIM805 : OR2B
      port map(A => \time_mem_wen_i_0[1]\, B => 
        time_mem_wen_i_0_0, Y => N_162);
    
    sFull_RNO_4 : OR2B
      port map(A => I_5_9, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[1]\);
    
    sFull_RNO_6 : OR2A
      port map(A => un1_waddr_vect_s, B => \time_mem_addr_w_1[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    sEmpty_RNO_3 : AX1E
      port map(A => un2_raddr_vect_s, B => I_9_10, C => 
        \Waddr_vect[2]_net_1\, Y => sEmpty_RNO_3_1);
    
    \Raddr_vect[2]\ : DFN1C0
      port map(D => Raddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Raddr_vect[2]_net_1\);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_1[0]\);
    
    sFull_RNO_5 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_9, C => 
        \Raddr_vect[2]_net_1\, Y => sFull_RNO_5_0);
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => \Waddr_vect[2]_net_1\, S
         => \time_mem_wen_i_0[1]\, Y => Waddr_vect_e2);
    
    un31_mem_addr_ren_I_8 : OR2B
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_1[5]\);
    
    sEmpty_RNO_4 : AX1E
      port map(A => un2_raddr_vect_s, B => I_5_10, C => 
        \time_mem_addr_w_1[1]\, Y => sEmpty_RNO_4_1);
    
    sFull_RNO_3 : XA1
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \un8_waddr_vect_s[3]\, C => time_ren(1), Y => 
        un5_sfull_s_2);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => sEmpty_RNO_3_1, B => sEmpty_RNO_4_1, C => 
        un7_sempty_s_0, Y => un7_sempty_s_3);
    
    \Waddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_w_1[0]\, B => 
        \time_mem_addr_w_1[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_n2_tz);
    
    un36_mem_addr_wen_I_5 : XOR2
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_1[3]\);
    
    \Raddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_r_1[0]\, B => 
        \time_mem_addr_r_1[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        Raddr_vect_n2_tz);
    
    sEmpty_RNO_7 : OR2A
      port map(A => un2_raddr_vect_s, B => \time_mem_addr_r_1[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Raddr_vect_RNO[2]\ : MX2A
      port map(A => Raddr_vect_n2, B => \Raddr_vect[2]_net_1\, S
         => \time_mem_ren_i_0[1]\, Y => Raddr_vect_e2);
    
    \Raddr_vect_RNIEJMC[3]\ : OR2B
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, Y => un2_raddr_vect_s);
    
    \Raddr_vect[0]\ : DFN1C0
      port map(D => Raddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_1[0]\);
    
    \sEmpty_RNI5EFO_0\ : OR2
      port map(A => \time_mem_ren_i_0[1]\, B => 
        \time_mem_addr_r_1[3]\, Y => sEmpty_RNI5EFO_0);
    
    \Raddr_vect_RNIHOG9[1]\ : OR3
      port map(A => \time_mem_addr_r_1[0]\, B => 
        \time_mem_addr_r_1[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        un2_raddr_vect_slt3);
    
    \Waddr_vect_RNINV58[2]\ : OR2A
      port map(A => \Waddr_vect[2]_net_1\, B => N_167, Y => 
        Waddr_vect_RNINV58(2));
    
    \Raddr_vect_RNI8J9L[2]\ : OR2A
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \time_mem_ren_i_0[1]\, Y => Raddr_vect_RNI8J9L(2));
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_r_1[1]\, B => 
        \time_mem_addr_r_1[0]\, Y => N_7);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_7_0, B => \Waddr_vect[2]_net_1\, Y => I_9_9);
    
    sFull_RNIC4G2 : OR2
      port map(A => time_wen(1), B => \sFull\, Y => 
        \time_mem_wen_i_0[1]\);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_4_0, B => \Raddr_vect[3]_net_1\, Y => 
        I_13_10);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_r_1[0]\, B => 
        \time_mem_addr_r_1[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        N_4_0);
    
    sEmpty_RNO_1 : XA1B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \un10_raddr_vect_s[3]\, C => time_ren(1), Y => 
        un7_sempty_s_2);
    
    sFull_RNO_1 : XA1
      port map(A => \un8_waddr_vect_s[1]\, B => 
        \time_mem_addr_r_1[1]\, C => sFull_RNO_5_0, Y => 
        un5_sfull_s_1);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_r_1[0]\, B => 
        \time_mem_addr_r_1[1]\, Y => I_5_10);
    
    \Waddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_w_1[0]\, B => 
        \time_mem_addr_w_1[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_15_0);
    
    sFull_RNO_7 : OR2B
      port map(A => I_13_9, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    \Raddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_r_1[0]\, B => 
        \time_mem_addr_r_1[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        Raddr_vect_7_0);
    
    \Raddr_vect_RNI6B9L[0]\ : OR2
      port map(A => \time_mem_ren_i_0[1]\, B => 
        \time_mem_addr_r_1[0]\, Y => N_70);
    
    \Waddr_vect_RNIMR58[1]\ : OR2
      port map(A => \time_mem_addr_w_1[1]\, B => N_167, Y => 
        N_146);
    
    \Waddr_vect_RNILN58[0]\ : OR2
      port map(A => \time_mem_addr_w_1[0]\, B => N_167, Y => 
        Waddr_vect_RNILN58(0));
    
    \Waddr_vect_RNO[3]\ : AXOI1
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, C => Waddr_vect_15_0, Y => 
        Waddr_vect_n3);
    
    un31_mem_addr_ren_I_16 : NOR2B
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \Raddr_vect[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    
    sFull_RNO_0 : NOR3C
      port map(A => un5_sfull_s_1, B => un5_sfull_s_0, C => 
        un5_sfull_s_2, Y => un5_sfull_s);
    
    sEmpty_RNO_6 : OR2B
      port map(A => I_13_10, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO_2\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \Waddr_vect_RNI2KMC[3]\ : OR2B
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, Y => un1_waddr_vect_s);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_1[1]\);
    
    sFull_RNO_2 : XA1B
      port map(A => \un8_waddr_vect_s[0]\, B => 
        \time_mem_addr_r_1[0]\, C => time_wen(1), Y => 
        un5_sfull_s_0);
    
    sEmpty_RNO_5 : XA1
      port map(A => \un10_raddr_vect_s[0]\, B => 
        \time_mem_addr_w_1[0]\, C => time_wen(1), Y => 
        un7_sempty_s_0);
    
    \Raddr_vect_RNO[3]\ : AXOI1
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, C => Raddr_vect_7_0, Y => 
        Raddr_vect_n3);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    sEmpty_RNICS3I : OR2
      port map(A => time_ren(1), B => \sEmpty\, Y => 
        \time_mem_ren_i_0[1]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ3 is

    port( ready_i_0          : out   std_logic_vector(3 to 3);
          data_mem_wen_i_0_0 : in    std_logic;
          data_ren           : in    std_logic_vector(3 to 3);
          data_wen           : in    std_logic_vector(3 to 3);
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic;
          N_128              : out   std_logic;
          N_152              : out   std_logic;
          N_136              : out   std_logic;
          N_68               : out   std_logic;
          N_144              : out   std_logic;
          N_166              : in    std_logic;
          N_160              : out   std_logic;
          N_76               : out   std_logic;
          N_60               : out   std_logic;
          N_52               : out   std_logic;
          N_86               : in    std_logic;
          N_44               : out   std_logic;
          N_1_i_1            : out   std_logic;
          N_1_i_1_i          : out   std_logic
        );

end lpp_waveform_fifo_ctrlZ3;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ3 is 

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_12, \data_mem_addr_w_3[1]\, \data_mem_addr_w_3[0]\, 
        N_4, \data_mem_addr_w_3[3]\, \DWACT_FINC_E[0]\, N_12_0, 
        \data_mem_addr_r_3[1]\, \data_mem_addr_r_3[0]\, N_4_0, 
        \data_mem_addr_r_3[3]\, \DWACT_FINC_E_0[0]\, 
        un7_sempty_s_4, un7_sempty_s_1, un7_sempty_s_0, 
        un7_sempty_s_2, \un10_raddr_vect_s[3]\, sEmpty_RNO_6_0, 
        \un10_raddr_vect_s[1]\, sEmpty_RNO_5_0, 
        \un10_raddr_vect_s[0]\, un5_sfull_s_4_2, 
        \un8_waddr_vect_s[3]\, \sFull_RNO_8\, un5_sfull_s_4_1, 
        \un8_waddr_vect_s[1]\, sFull_RNO_5_1, un5_sfull_s_4_0, 
        \un8_waddr_vect_s[0]\, ADD_7x7_fast_I23_Y_0_o2_0, N165_1, 
        \un174_ready0_1[4]\, N_11, ADD_5x5_fast_I11_Y_0, N80, 
        ADD_5x5_fast_I11_Y_i_a2_0, \data_mem_addr_w_3[2]\, 
        \data_mem_addr_r_3[2]\, \un189_ready0_1[4]\, 
        ADD_7x7_fast_I19_Y_i_o4_1_0, N_87, un1_waddr_vect_slto3_0, 
        un2_raddr_vect_slto3_0, I11_un1_Y, N81, N77, N98, N_12_1, 
        N_17, N_18, \un174_ready1[4]\, CO1_tz, un5_sfull_s_4, N_9, 
        Waddr_vect_n4, \data_mem_addr_w_3[4]\, Waddr_vect_14_0, 
        un1_waddr_vect_s, Waddr_vect_c2, Waddr_vect_n2, 
        Waddr_vect_c1, Waddr_vect_n3, N_105, \sFull_RNO_6\, 
        \sFull\, un1_sempty_s, \sEmpty\, sEmpty_RNO_8, I_5_11, 
        I_13_11, un2_raddr_vect_s, un2_raddr_vect_slto1, 
        \data_mem_addr_r_3[4]\, \un10_raddr_vect_s[2]\, 
        \un10_raddr_vect_s[4]\, \N_1_i_1\, \data_mem_wen_i_0[3]\, 
        N_75, N_24, N165, Waddr_vect_e2, Waddr_vect_e3, 
        Waddr_vect_e4, N111, N107, \un189_ready1_i[5]\, N_13, 
        N161, N_16_i, un191_ready, N_197_i, N_196_i, N_198, 
        \un189_ready1[4]\, \un189_ready0[4]\, un176_readylto4_i_0, 
        \un174_ready0[4]\, un183_ready, Waddr_vect_e0, 
        Waddr_vect_e1, Waddr_vect_n1_i, I_20_3, I_9_11, I_20_4, 
        I_13_12, I_9_12, I_5_12, sREN, N_9_0, N_13_0, N_12_2, 
        N_11_0, N_8, N_10, N_9_1, N_7, N_4_1, N_5, N_6, N_9_2, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    N_1_i_1 <= \N_1_i_1\;

    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \data_mem_addr_w_3[1]\, B => 
        \data_mem_addr_w_3[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_w_3[0]\, B => 
        \data_mem_addr_w_3[1]\, C => \data_mem_addr_w_3[2]\, Y
         => N_9_2);
    
    un189_ready_0_0_0_ADD_7x7_fast_I23_Y_0 : OR3A
      port map(A => N_75, B => N_24, C => 
        ADD_7x7_fast_I23_Y_0_o2_0, Y => N161);
    
    \ready_gen.un183_ready_0_I_9\ : AO1C
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \data_mem_addr_r_3[3]\, C => N_7, Y => N_12_2);
    
    un189_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4 : OR2B
      port map(A => N80, B => N165_1, Y => N165);
    
    \ready_gen.un183_ready_0_I_3\ : NOR2A
      port map(A => \data_mem_addr_r_3[0]\, B => 
        \data_mem_addr_w_3[0]\, Y => N_6);
    
    \Raddr_vect_RNIDKRC[4]\ : NOR2B
      port map(A => I_9_12, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[2]\);
    
    \Raddr_vect_RNI3FG82[0]\ : MX2C
      port map(A => N107, B => N161, S => \data_mem_addr_r_3[0]\, 
        Y => N_198);
    
    un189_ready_1_16_ADD_5x5_fast_I11_Y_0 : MIN3
      port map(A => \un174_ready0_1[4]\, B => N_11, C => N80, Y
         => ADD_5x5_fast_I11_Y_0);
    
    un189_ready_1_16_ADD_5x5_fast_I1_G0N : AO1C
      port map(A => \data_mem_addr_w_3[2]\, B => 
        \data_mem_addr_r_3[2]\, C => N_87, Y => N80);
    
    un8_raddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_r_3[0]\, B => 
        \data_mem_addr_r_3[1]\, C => \data_mem_addr_r_3[2]\, Y
         => \DWACT_FINC_E_0[0]\);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_w_3[1]\, B => 
        \data_mem_addr_w_3[0]\, Y => N_12);
    
    sEmpty_RNO : AO1A
      port map(A => data_ren(3), B => un7_sempty_s_4, C => 
        un1_sempty_s, Y => sEmpty_RNO_8);
    
    \Raddr_vect_RNIJBIK8[3]\ : OR2A
      port map(A => N_86, B => \data_mem_addr_r_3[3]\, Y => N_52);
    
    \ready_gen.un183_ready_0_I_1\ : OR2A
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \data_mem_addr_w_3[1]\, Y => N_4_1);
    
    \Raddr_vect[1]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sREN, Q => \data_mem_addr_r_3[1]\);
    
    \Waddr_vect[3]\ : DFN1C0
      port map(D => Waddr_vect_e3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_3[3]\);
    
    un189_ready_0_0_0_ADD_7x7_fast_I23_Y_0_a4_0 : NOR2A
      port map(A => N165, B => \un174_ready0_1[4]\, Y => N_24);
    
    \ready_gen.un183_ready_0_I_2\ : OR2A
      port map(A => \data_mem_addr_w_3[2]\, B => 
        \data_mem_addr_r_3[2]\, Y => N_5);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_12_0, B => \data_mem_addr_r_3[2]\, Y => 
        I_9_12);
    
    \Raddr_vect_RNIAG18[4]\ : AO1B
      port map(A => un2_raddr_vect_slto3_0, B => 
        un2_raddr_vect_slto1, C => \data_mem_addr_r_3[4]\, Y => 
        un2_raddr_vect_s);
    
    \Raddr_vect_RNISKHJ1[0]\ : MX2C
      port map(A => \un189_ready1[4]\, B => \un189_ready0[4]\, S
         => \data_mem_addr_r_3[0]\, Y => N_196_i);
    
    \Waddr_vect_RNO[4]\ : MX2A
      port map(A => Waddr_vect_n4, B => \data_mem_addr_w_3[4]\, S
         => \data_mem_wen_i_0[3]\, Y => Waddr_vect_e4);
    
    sEmpty : DFN1P0
      port map(D => sEmpty_RNO_8, CLK => HCLK_c, PRE => HRESETn_c, 
        Q => \sEmpty\);
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => \data_mem_wen_i_0[3]\, 
        C => \data_mem_addr_w_3[0]\, Y => Waddr_vect_e0);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_3[2]\);
    
    \ready_gen.un183_ready_0_I_6\ : OA1A
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \data_mem_addr_r_3[3]\, C => N_5, Y => N_9_1);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \data_mem_addr_w_3[1]\, 
        S => \data_mem_wen_i_0[3]\, Y => Waddr_vect_e1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un174_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0_0 : OA1A
      port map(A => \data_mem_addr_w_3[2]\, B => 
        \data_mem_addr_r_3[2]\, C => N_11, Y => 
        ADD_5x5_fast_I11_Y_i_a2_0);
    
    \Raddr_vect_RNIK03G[4]\ : NOR2B
      port map(A => I_20_4, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[4]\);
    
    \Waddr_vect_RNO_0[2]\ : XAI1A
      port map(A => \data_mem_addr_w_3[2]\, B => Waddr_vect_c1, C
         => un1_waddr_vect_s, Y => Waddr_vect_n2);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_w_3[0]\, B => 
        \data_mem_addr_w_3[1]\, Y => I_5_11);
    
    \Raddr_vect_RNIGVHK8[0]\ : OR2A
      port map(A => N_86, B => \data_mem_addr_r_3[0]\, Y => N_76);
    
    un174_ready_1_1_0_CO1_tz : AO18
      port map(A => N_105, B => \data_mem_addr_w_3[2]\, C => 
        \data_mem_addr_r_3[2]\, Y => CO1_tz);
    
    \Waddr_vect_RNIRR791[1]\ : OR3
      port map(A => N_166, B => data_mem_wen_i_0_0, C => 
        \data_mem_addr_w_3[1]\, Y => N_152);
    
    \ready_gen.un183_ready_0_I_7\ : AO1C
      port map(A => \data_mem_addr_w_3[2]\, B => 
        \data_mem_addr_r_3[2]\, C => N_4_1, Y => N_10);
    
    un189_ready_1_16_ADD_5x5_fast_I15_Y_0 : XOR2
      port map(A => N111, B => \un189_ready0_1[4]\, Y => 
        \un189_ready1[4]\);
    
    \Raddr_vect_RNIR7VE2[0]\ : MX2
      port map(A => \un189_ready1_i[5]\, B => N_16_i, S => 
        \data_mem_addr_r_3[0]\, Y => N_197_i);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sREN, Q => \data_mem_addr_r_3[3]\);
    
    sEmpty_RNO_2 : XA1A
      port map(A => \data_mem_addr_w_3[1]\, B => 
        \un10_raddr_vect_s[1]\, C => sEmpty_RNO_5_0, Y => 
        un7_sempty_s_1);
    
    \ready_gen.un183_ready_0_I_4\ : OR2A
      port map(A => \data_mem_addr_r_3[4]\, B => 
        \data_mem_addr_w_3[4]\, Y => N_7);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_9_2, B => \data_mem_addr_w_3[3]\, Y => 
        I_13_11);
    
    un174_ready_1_1_0_SUM2_0_0 : XOR2
      port map(A => N_11, B => \un174_ready0_1[4]\, Y => 
        \un189_ready0_1[4]\);
    
    \Waddr_vect_RNIBK63[0]\ : OR2B
      port map(A => \data_mem_addr_w_3[1]\, B => 
        \data_mem_addr_w_3[0]\, Y => Waddr_vect_c1);
    
    sFull_RNO : OA1
      port map(A => \sFull\, B => un5_sfull_s_4, C => data_ren(3), 
        Y => \sFull_RNO_6\);
    
    un189_ready_0_0_0_ADD_7x7_fast_I33_Y_0_i_x2 : AX1B
      port map(A => N_24, B => ADD_7x7_fast_I23_Y_0_o2_0, C => 
        N_75, Y => N_16_i);
    
    un189_ready_1_16_ADD_5x5_fast_I11_un1_Y : NOR3C
      port map(A => N81, B => N77, C => N98, Y => I11_un1_Y);
    
    un189_ready_0_0_0_ADD_7x7_fast_I32_Y_0 : XOR2
      port map(A => N165, B => \un189_ready0_1[4]\, Y => 
        \un189_ready0[4]\);
    
    \Raddr_vect_RNII7IK8[2]\ : OR2A
      port map(A => N_86, B => \data_mem_addr_r_3[2]\, Y => N_60);
    
    sFull_RNO_4 : OR2B
      port map(A => I_5_11, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[1]\);
    
    sFull_RNO_6 : OR2A
      port map(A => un1_waddr_vect_s, B => \data_mem_addr_w_3[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    sEmpty_RNO_3 : XA1A
      port map(A => \data_mem_addr_w_3[0]\, B => 
        \un10_raddr_vect_s[0]\, C => data_wen(3), Y => 
        un7_sempty_s_0);
    
    \Raddr_vect[2]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sREN, Q => \data_mem_addr_r_3[2]\);
    
    \Raddr_vect_RNIQB1B6[0]\ : AO1
      port map(A => N_197_i, B => N_196_i, C => N_198, Y => 
        un191_ready);
    
    un189_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1 : OR2B
      port map(A => ADD_7x7_fast_I19_Y_i_o4_1_0, B => N_9, Y => 
        N165_1);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_3[0]\);
    
    sFull_RNO_8 : AX1E
      port map(A => un1_waddr_vect_s, B => I_20_3, C => 
        \data_mem_addr_r_3[4]\, Y => \sFull_RNO_8\);
    
    un6_waddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \DWACT_FINC_E[0]\, Y => N_4);
    
    un174_ready_0_0_0_ADD_5x5_fast_I11_Y_i_o2 : OR2A
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \data_mem_addr_r_3[3]\, Y => N_11);
    
    sFull_RNO_5 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_11, C => 
        \data_mem_addr_r_3[2]\, Y => sFull_RNO_5_1);
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => \data_mem_addr_w_3[2]\, S
         => \data_mem_wen_i_0[3]\, Y => Waddr_vect_e2);
    
    \Raddr_vect_RNI5473[3]\ : NOR2
      port map(A => \data_mem_addr_r_3[3]\, B => 
        \data_mem_addr_r_3[2]\, Y => un2_raddr_vect_slto3_0);
    
    sEmpty_RNO_4 : XA1A
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \un10_raddr_vect_s[3]\, C => sEmpty_RNO_6_0, Y => 
        un7_sempty_s_2);
    
    \Waddr_vect_RNO_1[4]\ : OR2B
      port map(A => Waddr_vect_c2, B => \data_mem_addr_w_3[3]\, Y
         => Waddr_vect_14_0);
    
    sFull_RNO_3 : XA1
      port map(A => \data_mem_addr_r_3[3]\, B => 
        \un8_waddr_vect_s[3]\, C => \sFull_RNO_8\, Y => 
        un5_sfull_s_4_2);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => un7_sempty_s_1, B => un7_sempty_s_0, C => 
        un7_sempty_s_2, Y => un7_sempty_s_4);
    
    sEmpty_RNICNF32 : OR2
      port map(A => \sEmpty\, B => data_ren(3), Y => sREN);
    
    \ready_gen.un183_ready_0_I_11\ : OA1
      port map(A => N_13_0, B => N_12_2, C => N_11_0, Y => 
        un183_ready);
    
    \Raddr_vect_RNIAOK9[0]\ : NOR2A
      port map(A => un2_raddr_vect_s, B => \data_mem_addr_r_3[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    \Raddr_vect_RNIB48B[4]\ : NOR2B
      port map(A => I_5_12, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[1]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Raddr_vect_RNIDG73[4]\ : NOR2A
      port map(A => \data_mem_addr_r_3[4]\, B => 
        \data_mem_addr_w_3[4]\, Y => N_75);
    
    \Raddr_vect_RNIF2GJ8[0]\ : MX2
      port map(A => un176_readylto4_i_0, B => un191_ready, S => 
        un183_ready, Y => ready_i_0(3));
    
    un174_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3 : OR2A
      port map(A => N_9, B => \data_mem_addr_r_3[2]\, Y => N_17);
    
    \Raddr_vect[0]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sREN, Q => \data_mem_addr_r_3[0]\);
    
    un189_ready_1_16_ADD_5x5_fast_I2_P0N : OR2B
      port map(A => N_11, B => \un174_ready0_1[4]\, Y => N98);
    
    un174_ready_0_0_0_ADD_5x5_fast_I18_Y_0_1 : XNOR2
      port map(A => \data_mem_addr_w_3[4]\, B => 
        \data_mem_addr_r_3[4]\, Y => \un174_ready0_1[4]\);
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \data_mem_addr_r_3[0]\, Y => N_12_0);
    
    un189_ready_1_16_ADD_5x5_fast_I8_Y : AO1B
      port map(A => N81, B => N77, C => N80, Y => N111);
    
    un189_ready_1_16_ADD_5x5_fast_I0_CO1 : XA1B
      port map(A => \data_mem_addr_r_3[2]\, B => 
        \data_mem_addr_w_3[2]\, C => N_105, Y => N77);
    
    \Waddr_vect_RNI3H18[4]\ : AO1B
      port map(A => un1_waddr_vect_slto3_0, B => Waddr_vect_c1, C
         => \data_mem_addr_w_3[4]\, Y => un1_waddr_vect_s);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_12, B => \data_mem_addr_w_3[2]\, Y => 
        I_9_11);
    
    sFull_RNI4FGH1_0 : INV
      port map(A => \N_1_i_1\, Y => N_1_i_1_i);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_9_0, B => \data_mem_addr_r_3[3]\, Y => 
        I_13_12);
    
    un174_ready_0_0_0_ADD_5x5_fast_I18_Y_0 : AX1C
      port map(A => N_12_1, B => N_13, C => \un174_ready0_1[4]\, 
        Y => \un174_ready0[4]\);
    
    \Raddr_vect_RNI04FB1[0]\ : MX2C
      port map(A => \un174_ready1[4]\, B => \un174_ready0[4]\, S
         => \data_mem_addr_r_3[0]\, Y => un176_readylto4_i_0);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_r_3[0]\, B => 
        \data_mem_addr_r_3[1]\, C => \data_mem_addr_r_3[2]\, Y
         => N_9_0);
    
    un189_ready_1_16_ADD_5x5_fast_I10_Y : AO1B
      port map(A => N111, B => N98, C => N_75, Y => N107);
    
    \ready_gen.un183_ready_0_I_10\ : OA1A
      port map(A => N_8, B => N_10, C => N_9_1, Y => N_13_0);
    
    sEmpty_RNO_1 : NOR2B
      port map(A => \sEmpty\, B => data_wen(3), Y => un1_sempty_s);
    
    un8_raddr_vect_s_I_20 : XOR2
      port map(A => N_4_0, B => \data_mem_addr_r_3[4]\, Y => 
        I_20_4);
    
    \Raddr_vect_RNIB873[3]\ : XNOR2
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \data_mem_addr_r_3[3]\, Y => N_87);
    
    sFull_RNO_1 : XA1
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \un8_waddr_vect_s[1]\, C => sFull_RNO_5_1, Y => 
        un5_sfull_s_4_1);
    
    \Waddr_vect_RNIT3891[3]\ : OR3
      port map(A => N_166, B => data_mem_wen_i_0_0, C => 
        \data_mem_addr_w_3[3]\, Y => N_136);
    
    \Waddr_vect_RNII4Q4[2]\ : NOR2A
      port map(A => \data_mem_addr_w_3[2]\, B => Waddr_vect_c1, Y
         => Waddr_vect_c2);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_r_3[0]\, B => 
        \data_mem_addr_r_3[1]\, Y => I_5_12);
    
    un189_ready_0_0_0_ADD_7x7_fast_I23_Y_0_o2_0 : AOI1
      port map(A => N165_1, B => \un174_ready0_1[4]\, C => N_11, 
        Y => ADD_7x7_fast_I23_Y_0_o2_0);
    
    un174_ready_0_0_0_ADD_5x5_fast_I9_Y_i_o2 : AO13
      port map(A => \data_mem_addr_w_3[1]\, B => 
        \data_mem_addr_w_3[0]\, C => \data_mem_addr_r_3[1]\, Y
         => N_9);
    
    \Waddr_vect_RNIF473[3]\ : NOR2
      port map(A => \data_mem_addr_w_3[3]\, B => 
        \data_mem_addr_w_3[2]\, Y => un1_waddr_vect_slto3_0);
    
    un189_ready_1_16_ADD_5x5_fast_I16_Y_0 : AX1B
      port map(A => I11_un1_Y, B => ADD_5x5_fast_I11_Y_0, C => 
        N_75, Y => \un189_ready1_i[5]\);
    
    \Raddr_vect_RNI7O63[1]\ : NOR2A
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \data_mem_addr_w_3[1]\, Y => N_105);
    
    \Raddr_vect_RNI1K63[1]\ : OR2B
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \data_mem_addr_r_3[0]\, Y => un2_raddr_vect_slto1);
    
    \Waddr_vect_RNO_0[3]\ : XAI1
      port map(A => \data_mem_addr_w_3[3]\, B => Waddr_vect_c2, C
         => un1_waddr_vect_s, Y => Waddr_vect_n3);
    
    \Waddr_vect[4]\ : DFN1C0
      port map(D => Waddr_vect_e4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_3[4]\);
    
    sFull_RNO_7 : OR2B
      port map(A => I_13_11, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    \Waddr_vect_RNIU7891[4]\ : OR3
      port map(A => N_166, B => data_mem_wen_i_0_0, C => 
        \data_mem_addr_w_3[4]\, Y => N_128);
    
    \Waddr_vect_RNIQN791[0]\ : OR3
      port map(A => N_166, B => data_mem_wen_i_0_0, C => 
        \data_mem_addr_w_3[0]\, Y => N_160);
    
    un174_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3_0 : OR2B
      port map(A => N_9, B => \data_mem_addr_w_3[2]\, Y => N_18);
    
    sFull_RNI4FGH1 : OR3A
      port map(A => \data_mem_wen_i_0[3]\, B => N_166, C => 
        data_mem_wen_i_0_0, Y => \N_1_i_1\);
    
    \Waddr_vect_RNO[3]\ : MX2A
      port map(A => Waddr_vect_n3, B => \data_mem_addr_w_3[3]\, S
         => \data_mem_wen_i_0[3]\, Y => Waddr_vect_e3);
    
    un189_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1_0 : AXOI5
      port map(A => N_87, B => \data_mem_addr_r_3[2]\, C => 
        \data_mem_addr_w_3[2]\, Y => ADD_7x7_fast_I19_Y_i_o4_1_0);
    
    un174_ready_1_1_0_SUM2_0 : AX1E
      port map(A => N_87, B => CO1_tz, C => \un189_ready0_1[4]\, 
        Y => \un174_ready1[4]\);
    
    un174_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2 : OR3C
      port map(A => N_17, B => ADD_5x5_fast_I11_Y_i_a2_0, C => 
        N_18, Y => N_12_1);
    
    sFull_RNO_0 : NOR3C
      port map(A => un5_sfull_s_4_1, B => un5_sfull_s_4_0, C => 
        un5_sfull_s_4_2, Y => un5_sfull_s_4);
    
    sEmpty_RNO_6 : XNOR2
      port map(A => \un10_raddr_vect_s[4]\, B => 
        \data_mem_addr_w_3[4]\, Y => sEmpty_RNO_6_0);
    
    \Waddr_vect_RNISV791[2]\ : OR3
      port map(A => N_166, B => data_mem_wen_i_0_0, C => 
        \data_mem_addr_w_3[2]\, Y => N_144);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO_6\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \Raddr_vect_RNIG8FE[4]\ : NOR2B
      port map(A => I_13_12, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    un6_waddr_vect_s_I_20 : XOR2
      port map(A => N_4, B => \data_mem_addr_w_3[4]\, Y => I_20_3);
    
    \ready_gen.un183_ready_0_I_8\ : OR2A
      port map(A => \data_mem_addr_w_3[4]\, B => 
        \data_mem_addr_r_3[4]\, Y => N_11_0);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_3[1]\);
    
    \ready_gen.un183_ready_0_I_5\ : AO1C
      port map(A => \data_mem_addr_r_3[1]\, B => 
        \data_mem_addr_w_3[1]\, C => N_6, Y => N_8);
    
    \Raddr_vect[4]\ : DFN1E0C0
      port map(D => \un10_raddr_vect_s[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => sREN, Q => \data_mem_addr_r_3[4]\);
    
    sFull_RNO_2 : XA1B
      port map(A => \data_mem_addr_r_3[0]\, B => 
        \un8_waddr_vect_s[0]\, C => data_wen(3), Y => 
        un5_sfull_s_4_0);
    
    un8_raddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_r_3[3]\, B => 
        \DWACT_FINC_E_0[0]\, Y => N_4_0);
    
    un174_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0 : OR2A
      port map(A => \data_mem_addr_r_3[3]\, B => 
        \data_mem_addr_w_3[3]\, Y => N_13);
    
    sEmpty_RNO_5 : XNOR2
      port map(A => \un10_raddr_vect_s[2]\, B => 
        \data_mem_addr_w_3[2]\, Y => sEmpty_RNO_5_0);
    
    \Raddr_vect_RNIKFIK8[4]\ : OR2A
      port map(A => N_86, B => \data_mem_addr_r_3[4]\, Y => N_44);
    
    \Raddr_vect_RNIH3IK8[1]\ : OR2A
      port map(A => N_86, B => \data_mem_addr_r_3[1]\, Y => N_68);
    
    sFull_RNIFVR9 : OR2
      port map(A => \sFull\, B => data_wen(3), Y => 
        \data_mem_wen_i_0[3]\);
    
    \Waddr_vect_RNO_0[4]\ : XAI1A
      port map(A => \data_mem_addr_w_3[4]\, B => Waddr_vect_14_0, 
        C => un1_waddr_vect_s, Y => Waddr_vect_n4);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un6_waddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_w_3[0]\, B => 
        \data_mem_addr_w_3[1]\, C => \data_mem_addr_w_3[2]\, Y
         => \DWACT_FINC_E[0]\);
    
    un189_ready_1_16_ADD_5x5_fast_I1_P0N : OR3A
      port map(A => \data_mem_addr_r_3[2]\, B => 
        \data_mem_addr_w_3[2]\, C => N_87, Y => N81);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ0 is

    port( ready_i_0                   : out   std_logic_vector(0 to 0);
          data_ren                    : in    std_logic_vector(0 to 0);
          data_addr_w_0_iv_i_1        : in    std_logic_vector(5 to 5);
          data_addr_r_1_iv_i_s_1      : in    std_logic_vector(6 to 6);
          data_addr_r_1_iv_i_a9_1_1   : in    std_logic_vector(6 to 6);
          data_mem_ren_i_0            : out   std_logic_vector(0 to 0);
          data_mem_wen_i_0_1          : in    std_logic;
          data_addr_w_1_iv_i_a2_1_1_0 : out   std_logic_vector(6 to 6);
          data_addr_w_iv_i_2          : in    std_logic_vector(4 downto 0);
          data_addr_w_iv_i_4          : out   std_logic_vector(4 downto 0);
          data_wen                    : in    std_logic_vector(0 to 0);
          data_addr_r_iv_i_0          : in    std_logic_vector(4 downto 0);
          data_addr_r_iv_i_1          : in    std_logic_vector(4 downto 0);
          data_addr_r_iv_i_3          : out   std_logic_vector(4 downto 0);
          HRESETn_c                   : in    std_logic;
          HCLK_c                      : in    std_logic;
          N_165                       : out   std_logic;
          N_120_i                     : in    std_logic;
          sFull_RNIHL443              : out   std_logic;
          sEmpty_RNILSD08             : out   std_logic;
          N_124                       : in    std_logic;
          N_164                       : in    std_logic;
          N_158                       : in    std_logic;
          N_142                       : in    std_logic;
          N_134                       : in    std_logic;
          N_126                       : in    std_logic;
          N_150                       : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ0;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ0 is 

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXO5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_12, \data_mem_addr_w_0[1]\, \data_mem_addr_w_0[0]\, 
        N_4, \data_mem_addr_w_0[3]\, \DWACT_FINC_E[0]\, N_12_0, 
        \data_mem_addr_r_0[1]\, \data_mem_addr_r_0[0]\, N_4_0, 
        \data_mem_addr_r_0[3]\, \DWACT_FINC_E_0[0]\, N_65, N_41, 
        N_49, N_57, N_73, un7_sempty_s_4, un7_sempty_s_1, 
        un7_sempty_s_0, un7_sempty_s_2, \un10_raddr_vect_s[3]\, 
        sEmpty_RNO_6_1, \un10_raddr_vect_s[1]\, sEmpty_RNO_5_1, 
        \un10_raddr_vect_s[0]\, N_149, N_125, N_133, N_141, N_157, 
        un5_sfull_s_4_2, \un8_waddr_vect_s[3]\, sFull_RNO_8_1, 
        un5_sfull_s_4_1, \un8_waddr_vect_s[1]\, sFull_RNO_5_3, 
        un5_sfull_s_4_0, \un8_waddr_vect_s[0]\, 
        \data_addr_w_0_iv_i_3[5]\, \data_mem_wen_i_0[0]\, 
        ADD_7x7_fast_I23_Y_0_o2_0, N165_1, N_89_i, N_109, 
        ADD_5x5_fast_I11_Y_0, N80, ADD_5x5_fast_I11_Y_i_a2_0, 
        \data_mem_addr_r_0[2]\, \data_mem_addr_w_0[2]\, SUM2_0_0, 
        ADD_7x7_fast_I19_Y_i_o4_1_0, N_87, un1_waddr_vect_slto3_0, 
        un2_raddr_vect_slto3_0, I11_un1_Y, N81, N77, N98, 
        \un3_ready1[4]\, CO1_tz, N_12_1, N_17, N_18, 
        un5_sfull_s_4, ADD_5x5_fast_I9_Y_i_o2_0, Waddr_vect_c1, 
        Waddr_vect_n4, \data_mem_addr_w_0[4]\, Waddr_vect_14_0, 
        un1_waddr_vect_s, Waddr_vect_c2, \sFull_RNO_7\, \sFull\, 
        Waddr_vect_n2, Waddr_vect_n3, N_84_1, 
        \data_mem_ren_i_0[0]\, \sEmpty\, un2_raddr_vect_s, I_5_14, 
        \un10_raddr_vect_s[2]\, I_9_14, I_13_14, 
        \un10_raddr_vect_s[4]\, I_20_6, un2_raddr_vect_slto1, 
        \data_mem_addr_r_0[4]\, I_9_13, ADD_5x5_fast_I8_un1_Y, 
        sEmpty_RNO_9, un1_sempty_s, N_75, Waddr_vect_e0, 
        Waddr_vect_e1, Waddr_vect_n1_i, Waddr_vect_e2, 
        Waddr_vect_e3, Waddr_vect_e4, \un18_ready1[4]\, 
        \un18_ready0_1[4]\, \un3_ready0[4]\, N_6, 
        \un18_ready0[4]\, un5_readylto4, un20_ready, un12_ready, 
        N_198, N107, N161, N_197, \un18_ready1[5]\, N_16_i_i_0, 
        N_196, N_24, N_13, I_20_5, I_13_13, I_5_13, N_9, N_13_0, 
        N_12_2, N_11, N_8, N_10, N_9_0, N_7, N_4_1, N_5, N_6_0, 
        N_9_1, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    data_mem_ren_i_0(0) <= \data_mem_ren_i_0[0]\;

    un3_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0_0 : AO1A
      port map(A => \data_mem_addr_r_0[2]\, B => 
        \data_mem_addr_w_0[2]\, C => N_109, Y => 
        ADD_5x5_fast_I11_Y_i_a2_0);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO_7\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \Waddr_vect_RNO[0]\ : AXOI5
      port map(A => un1_waddr_vect_s, B => \data_mem_wen_i_0[0]\, 
        C => \data_mem_addr_w_0[0]\, Y => Waddr_vect_e0);
    
    un3_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2_0 : OR2A
      port map(A => \data_mem_addr_r_0[3]\, B => 
        \data_mem_addr_w_0[3]\, Y => N_13);
    
    sFull_RNO_8 : AX1E
      port map(A => un1_waddr_vect_s, B => I_20_5, C => 
        \data_mem_addr_r_0[4]\, Y => sFull_RNO_8_1);
    
    \Waddr_vect_RNI11GL[2]\ : OR3A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => 
        \data_mem_addr_w_0[2]\, Y => N_141);
    
    \Waddr_vect_RNIC9KQ2[2]\ : NOR3C
      port map(A => N_141, B => data_addr_w_iv_i_2(2), C => N_142, 
        Y => data_addr_w_iv_i_4(2));
    
    sFull_RNO_6 : OR2A
      port map(A => un1_waddr_vect_s, B => \data_mem_addr_w_0[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    \Raddr_vect_RNI73352[1]\ : OR2A
      port map(A => \data_mem_ren_i_0[0]\, B => 
        \data_mem_addr_r_0[1]\, Y => N_65);
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_0[0]\);
    
    \Waddr_vect_RNO[3]\ : MX2B
      port map(A => \data_mem_addr_w_0[3]\, B => Waddr_vect_n3, S
         => \data_mem_wen_i_0[0]\, Y => Waddr_vect_e3);
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \data_mem_addr_r_0[0]\, Y => N_12_0);
    
    un18_ready_0_0_0_ADD_7x7_fast_I23_Y_0_a4_0 : AO1D
      port map(A => N80, B => N165_1, C => N_89_i, Y => N_24);
    
    \Waddr_vect_RNIKG18[4]\ : AO1B
      port map(A => un1_waddr_vect_slto3_0, B => Waddr_vect_c1, C
         => \data_mem_addr_w_0[4]\, Y => un1_waddr_vect_s);
    
    \Raddr_vect_RNILJRC[4]\ : NOR2B
      port map(A => I_9_14, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[2]\);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_w_0[0]\, B => 
        \data_mem_addr_w_0[1]\, Y => I_5_13);
    
    \ready_gen.un12_ready_0_I_10\ : OA1A
      port map(A => N_8, B => N_10, C => N_9_0, Y => N_13_0);
    
    \Raddr_vect_RNI5873[3]\ : XNOR2
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \data_mem_addr_r_0[3]\, Y => N_87);
    
    \Raddr_vect_RNIV373[3]\ : NOR2
      port map(A => \data_mem_addr_r_0[3]\, B => 
        \data_mem_addr_r_0[2]\, Y => un2_raddr_vect_slto3_0);
    
    \sFull_RNIHL443\ : NOR3C
      port map(A => data_addr_w_0_iv_i_1(5), B => N_120_i, C => 
        \data_addr_w_0_iv_i_3[5]\, Y => sFull_RNIHL443);
    
    \Raddr_vect_RNI87352[2]\ : OR2A
      port map(A => \data_mem_ren_i_0[0]\, B => 
        \data_mem_addr_r_0[2]\, Y => N_57);
    
    un18_ready_1_16_ADD_5x5_fast_I10_Y : OR3A
      port map(A => N_75, B => ADD_5x5_fast_I8_un1_Y, C => N80, Y
         => N107);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => un7_sempty_s_1, B => un7_sempty_s_0, C => 
        un7_sempty_s_2, Y => un7_sempty_s_4);
    
    \ready_gen.un12_ready_0_I_11\ : OA1
      port map(A => N_13_0, B => N_12_2, C => N_11, Y => 
        un12_ready);
    
    un18_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1_0 : AXO5
      port map(A => N_87, B => \data_mem_addr_r_0[2]\, C => 
        \data_mem_addr_w_0[2]\, Y => ADD_7x7_fast_I19_Y_i_o4_1_0);
    
    un18_ready_0_0_0_ADD_7x7_fast_I23_Y_0_o2_0 : AO1C
      port map(A => N165_1, B => N_89_i, C => N_109, Y => 
        ADD_7x7_fast_I23_Y_0_o2_0);
    
    \Waddr_vect_RNI94Q4[2]\ : NOR2A
      port map(A => \data_mem_addr_w_0[2]\, B => Waddr_vect_c1, Y
         => Waddr_vect_c2);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_r_0[0]\, B => 
        \data_mem_addr_r_0[1]\, C => \data_mem_addr_r_0[2]\, Y
         => N_9);
    
    un18_ready_1_16_ADD_5x5_fast_I11_Y_0 : AO18
      port map(A => N80, B => N_89_i, C => N_109, Y => 
        ADD_5x5_fast_I11_Y_0);
    
    \Waddr_vect_RNO[4]\ : MX2B
      port map(A => \data_mem_addr_w_0[4]\, B => Waddr_vect_n4, S
         => \data_mem_wen_i_0[0]\, Y => Waddr_vect_e4);
    
    un3_ready_1_1_0_SUM2_0 : AX1C
      port map(A => N_87, B => CO1_tz, C => SUM2_0_0, Y => 
        \un3_ready1[4]\);
    
    \Waddr_vect_RNI5K63[0]\ : OR2B
      port map(A => \data_mem_addr_w_0[1]\, B => 
        \data_mem_addr_w_0[0]\, Y => Waddr_vect_c1);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_0[1]\);
    
    \ready_gen.un12_ready_0_I_9\ : AO1C
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \data_mem_addr_r_0[3]\, C => N_7, Y => N_12_2);
    
    sFull_RNO_7 : OR2B
      port map(A => I_13_13, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_9_1, B => \data_mem_addr_w_0[3]\, Y => 
        I_13_13);
    
    GND_i : GND
      port map(Y => \GND\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \ready_gen.un12_ready_0_I_2\ : OR2A
      port map(A => \data_mem_addr_w_0[2]\, B => 
        \data_mem_addr_r_0[2]\, Y => N_5);
    
    \Waddr_vect_RNI0TFL[1]\ : OR3A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => 
        \data_mem_addr_w_0[1]\, Y => N_149);
    
    sFull_RNITGSJ : NOR2
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, Y => N_165);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \data_mem_addr_w_0[0]\, B => 
        \data_mem_addr_w_0[1]\, C => \data_mem_addr_w_0[2]\, Y
         => N_9_1);
    
    un18_ready_1_16_ADD_5x5_fast_I16_Y_0 : AX1E
      port map(A => I11_un1_Y, B => ADD_5x5_fast_I11_Y_0, C => 
        N_75, Y => \un18_ready1[5]\);
    
    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \data_mem_addr_w_0[1]\, B => 
        \data_mem_addr_w_0[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    \Raddr_vect_RNIMV2G[4]\ : NOR2B
      port map(A => I_20_6, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[4]\);
    
    \Raddr_vect[2]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[0]\, Q => 
        \data_mem_addr_r_0[2]\);
    
    \Raddr_vect_RNI48175[4]\ : NOR3C
      port map(A => data_addr_r_iv_i_1(4), B => 
        data_addr_r_iv_i_0(4), C => N_41, Y => 
        data_addr_r_iv_i_3(4));
    
    sFull_RNIKUNJ : NOR2A
      port map(A => data_mem_wen_i_0_1, B => 
        \data_mem_wen_i_0[0]\, Y => 
        data_addr_w_1_iv_i_a2_1_1_0(6));
    
    \Raddr_vect_RNI6V252[0]\ : OR2A
      port map(A => \data_mem_ren_i_0[0]\, B => 
        \data_mem_addr_r_0[0]\, Y => N_73);
    
    sFull_RNI9VR9 : NOR2
      port map(A => \sFull\, B => data_wen(0), Y => 
        \data_mem_wen_i_0[0]\);
    
    un18_ready_1_16_ADD_5x5_fast_I1_G0N : OA1A
      port map(A => \data_mem_addr_r_0[2]\, B => 
        \data_mem_addr_w_0[2]\, C => N_87, Y => N80);
    
    \ready_gen.un12_ready_0_I_7\ : AO1C
      port map(A => \data_mem_addr_w_0[2]\, B => 
        \data_mem_addr_r_0[2]\, C => N_4_1, Y => N_10);
    
    \Waddr_vect_RNO_0[4]\ : XAI1A
      port map(A => \data_mem_addr_w_0[4]\, B => Waddr_vect_14_0, 
        C => un1_waddr_vect_s, Y => Waddr_vect_n4);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un3_ready_0_0_0_ADD_5x5_fast_I11_Y_i : OR2B
      port map(A => N_13, B => N_12_1, Y => N_6);
    
    un18_ready_1_16_ADD_5x5_fast_I2_P0N : OR2A
      port map(A => N_89_i, B => N_109, Y => N98);
    
    sEmpty_RNO : AO1A
      port map(A => data_ren(0), B => un7_sempty_s_4, C => 
        un1_sempty_s, Y => sEmpty_RNO_9);
    
    \Raddr_vect_RNIONK9[0]\ : NOR2A
      port map(A => un2_raddr_vect_s, B => \data_mem_addr_r_0[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    \Raddr_vect_RNI6QHR1[0]\ : MX2C
      port map(A => N107, B => N161, S => \data_mem_addr_r_0[0]\, 
        Y => N_198);
    
    \Waddr_vect[3]\ : DFN1C0
      port map(D => Waddr_vect_e3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_0[3]\);
    
    un3_ready_1_1_0_CO1_tz : AO18
      port map(A => N_84_1, B => \data_mem_addr_w_0[2]\, C => 
        \data_mem_addr_r_0[2]\, Y => CO1_tz);
    
    un3_ready_0_0_0_ADD_5x5_fast_I9_Y_i_o2_0 : AO1D
      port map(A => \data_mem_addr_w_0[1]\, B => 
        \data_mem_addr_w_0[0]\, C => \data_mem_addr_r_0[1]\, Y
         => ADD_5x5_fast_I9_Y_i_o2_0);
    
    un18_ready_1_16_ADD_5x5_fast_I8_un1_Y : NOR2B
      port map(A => N81, B => N77, Y => ADD_5x5_fast_I8_un1_Y);
    
    un18_ready_1_16_ADD_5x5_fast_I15_Y_0 : AX1D
      port map(A => ADD_5x5_fast_I8_un1_Y, B => N80, C => 
        \un18_ready0_1[4]\, Y => \un18_ready1[4]\);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \data_mem_addr_w_0[1]\, B => 
        \data_mem_addr_w_0[0]\, Y => N_12);
    
    sEmpty_RNO_3 : XA1A
      port map(A => \data_mem_addr_w_0[0]\, B => 
        \un10_raddr_vect_s[0]\, C => data_wen(0), Y => 
        un7_sempty_s_0);
    
    \sEmpty_RNILSD08\ : AO1C
      port map(A => \data_mem_ren_i_0[0]\, B => 
        data_addr_r_1_iv_i_a9_1_1(6), C => 
        data_addr_r_1_iv_i_s_1(6), Y => sEmpty_RNILSD08);
    
    \Raddr_vect_RNIRF18[4]\ : AO1B
      port map(A => un2_raddr_vect_slto3_0, B => 
        un2_raddr_vect_slto1, C => \data_mem_addr_r_0[4]\, Y => 
        un2_raddr_vect_s);
    
    \Raddr_vect_RNIPBM76[0]\ : AOI1
      port map(A => N_197, B => N_196, C => N_198, Y => 
        un20_ready);
    
    un6_waddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \DWACT_FINC_E[0]\, Y => N_4);
    
    \Waddr_vect_RNI39GL[4]\ : OR3A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => 
        \data_mem_addr_w_0[4]\, Y => N_125);
    
    un3_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3_0 : AOI1B
      port map(A => ADD_5x5_fast_I9_Y_i_o2_0, B => Waddr_vect_c1, 
        C => \data_mem_addr_w_0[2]\, Y => N_18);
    
    \Waddr_vect[4]\ : DFN1C0
      port map(D => Waddr_vect_e4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_0[4]\);
    
    sFull_RNO : OA1
      port map(A => \sFull\, B => un5_sfull_s_4, C => data_ren(0), 
        Y => \sFull_RNO_7\);
    
    sFull_RNO_2 : XA1B
      port map(A => \data_mem_addr_r_0[0]\, B => 
        \un8_waddr_vect_s[0]\, C => data_wen(0), Y => 
        un5_sfull_s_4_0);
    
    un3_ready_0_0_0_ADD_5x5_fast_I11_Y_i_a2 : OR3
      port map(A => N_17, B => ADD_5x5_fast_I11_Y_i_a2_0, C => 
        N_18, Y => N_12_1);
    
    \Waddr_vect_RNO_0[2]\ : XAI1A
      port map(A => \data_mem_addr_w_0[2]\, B => Waddr_vect_c1, C
         => un1_waddr_vect_s, Y => Waddr_vect_n2);
    
    \Raddr_vect_RNIRJ63[1]\ : OR2B
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \data_mem_addr_r_0[0]\, Y => un2_raddr_vect_slto1);
    
    \Waddr_vect_RNIQ5C73[4]\ : NOR3C
      port map(A => N_125, B => data_addr_w_iv_i_2(4), C => N_126, 
        Y => data_addr_w_iv_i_4(4));
    
    \Raddr_vect[0]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[0]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[0]\, Q => 
        \data_mem_addr_r_0[0]\);
    
    \Waddr_vect_RNIQL7S2[3]\ : NOR3C
      port map(A => N_133, B => data_addr_w_iv_i_2(3), C => N_134, 
        Y => data_addr_w_iv_i_4(3));
    
    \Raddr_vect_RNI16OM1[0]\ : MX2C
      port map(A => \un18_ready1[4]\, B => \un18_ready0[4]\, S
         => \data_mem_addr_r_0[0]\, Y => N_196);
    
    \Waddr_vect_RNO_0[3]\ : XAI1
      port map(A => \data_mem_addr_w_0[3]\, B => Waddr_vect_c2, C
         => un1_waddr_vect_s, Y => Waddr_vect_n3);
    
    \Raddr_vect_RNIIBCL2[0]\ : MX2C
      port map(A => \un18_ready1[5]\, B => N_16_i_i_0, S => 
        \data_mem_addr_r_0[0]\, Y => N_197);
    
    \Raddr_vect_RNIL7FE[4]\ : NOR2B
      port map(A => I_13_14, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    \Raddr_vect_RNI5873_0[3]\ : NOR2A
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \data_mem_addr_r_0[3]\, Y => N_109);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_12_0, B => \data_mem_addr_r_0[2]\, Y => 
        I_9_14);
    
    un18_ready_0_0_0_ADD_7x7_fast_I33_Y_0_i_x2 : AX1E
      port map(A => N_24, B => ADD_7x7_fast_I23_Y_0_o2_0, C => 
        N_75, Y => N_16_i_i_0);
    
    un18_ready_1_16_ADD_5x5_fast_I1_P0N : OR3A
      port map(A => \data_mem_addr_r_0[2]\, B => 
        \data_mem_addr_w_0[2]\, C => N_87, Y => N81);
    
    sFull_RNO_3 : XA1
      port map(A => \data_mem_addr_r_0[3]\, B => 
        \un8_waddr_vect_s[3]\, C => sFull_RNO_8_1, Y => 
        un5_sfull_s_4_2);
    
    sEmpty_RNI9NF32 : NOR2
      port map(A => \sEmpty\, B => data_ren(0), Y => 
        \data_mem_ren_i_0[0]\);
    
    \ready_gen.un12_ready_0_I_6\ : OA1A
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \data_mem_addr_r_0[3]\, C => N_5, Y => N_9_0);
    
    un8_raddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_r_0[0]\, B => 
        \data_mem_addr_r_0[1]\, C => \data_mem_addr_r_0[2]\, Y
         => \DWACT_FINC_E_0[0]\);
    
    \Waddr_vect_RNO_1[4]\ : OR2B
      port map(A => Waddr_vect_c2, B => \data_mem_addr_w_0[3]\, Y
         => Waddr_vect_14_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un18_ready_0_0_0_ADD_7x7_fast_I23_Y_0 : OR2A
      port map(A => N_75, B => \un3_ready0[4]\, Y => N161);
    
    \Raddr_vect_RNI34175[3]\ : NOR3C
      port map(A => data_addr_r_iv_i_1(3), B => 
        data_addr_r_iv_i_0(3), C => N_49, Y => 
        data_addr_r_iv_i_3(3));
    
    un6_waddr_vect_s_I_20 : XOR2
      port map(A => N_4, B => \data_mem_addr_w_0[4]\, Y => I_20_5);
    
    \Raddr_vect[1]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[1]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[0]\, Q => 
        \data_mem_addr_r_0[1]\);
    
    sEmpty_RNO_6 : XNOR2
      port map(A => \un10_raddr_vect_s[4]\, B => 
        \data_mem_addr_w_0[4]\, Y => sEmpty_RNO_6_1);
    
    sFull_RNIOK841 : OA1A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => N_124, 
        Y => \data_addr_w_0_iv_i_3[5]\);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_9, B => \data_mem_addr_r_0[3]\, Y => 
        I_13_14);
    
    \Waddr_vect_RNO[2]\ : MX2B
      port map(A => \data_mem_addr_w_0[2]\, B => Waddr_vect_n2, S
         => \data_mem_wen_i_0[0]\, Y => Waddr_vect_e2);
    
    sFull_RNO_0 : NOR3C
      port map(A => un5_sfull_s_4_1, B => un5_sfull_s_4_0, C => 
        un5_sfull_s_4_2, Y => un5_sfull_s_4);
    
    \Raddr_vect_RNIAF352[4]\ : OR2A
      port map(A => \data_mem_ren_i_0[0]\, B => 
        \data_mem_addr_r_0[4]\, Y => N_41);
    
    sEmpty_RNO_2 : XA1A
      port map(A => \data_mem_addr_w_0[1]\, B => 
        \un10_raddr_vect_s[1]\, C => sEmpty_RNO_5_1, Y => 
        un7_sempty_s_1);
    
    \Raddr_vect_RNIP9SH1[0]\ : MX2
      port map(A => \un3_ready1[4]\, B => \un3_ready0[4]\, S => 
        \data_mem_addr_r_0[0]\, Y => un5_readylto4);
    
    \Raddr_vect_RNI1O63[1]\ : NOR2A
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \data_mem_addr_w_0[1]\, Y => N_84_1);
    
    sEmpty_RNO_4 : XA1A
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \un10_raddr_vect_s[3]\, C => sEmpty_RNO_6_1, Y => 
        un7_sempty_s_2);
    
    sFull_RNO_5 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_13, C => 
        \data_mem_addr_r_0[2]\, Y => sFull_RNO_5_3);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \data_mem_addr_r_0[0]\, B => 
        \data_mem_addr_r_0[1]\, Y => I_5_14);
    
    un18_ready_0_0_0_ADD_7x7_fast_I19_Y_i_o4_1 : AOI1
      port map(A => ADD_5x5_fast_I9_Y_i_o2_0, B => Waddr_vect_c1, 
        C => ADD_7x7_fast_I19_Y_i_o4_1_0, Y => N165_1);
    
    \ready_gen.un12_ready_0_I_8\ : OR2A
      port map(A => \data_mem_addr_w_0[4]\, B => 
        \data_mem_addr_r_0[4]\, Y => N_11);
    
    \Raddr_vect_RNIH6IM8[0]\ : MX2
      port map(A => un5_readylto4, B => un20_ready, S => 
        un12_ready, Y => ready_i_0(0));
    
    \Waddr_vect_RNI25GL[3]\ : OR3A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => 
        \data_mem_addr_w_0[3]\, Y => N_133);
    
    sEmpty : DFN1P0
      port map(D => sEmpty_RNO_9, CLK => HCLK_c, PRE => HRESETn_c, 
        Q => \sEmpty\);
    
    \Waddr_vect_RNO[1]\ : MX2B
      port map(A => \data_mem_addr_w_0[1]\, B => Waddr_vect_n1_i, 
        S => \data_mem_wen_i_0[0]\, Y => Waddr_vect_e1);
    
    un18_ready_0_0_0_ADD_7x7_fast_I32_Y_0_1 : XNOR2
      port map(A => N_109, B => N_89_i, Y => \un18_ready0_1[4]\);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_mem_addr_w_0[2]\);
    
    \Waddr_vect_RNI58KI2[0]\ : NOR3C
      port map(A => N_157, B => data_addr_w_iv_i_2(0), C => N_158, 
        Y => data_addr_w_iv_i_4(0));
    
    \Raddr_vect_RNI2C8Q4[0]\ : NOR3C
      port map(A => data_addr_r_iv_i_1(0), B => 
        data_addr_r_iv_i_0(0), C => N_73, Y => 
        data_addr_r_iv_i_3(0));
    
    un18_ready_0_0_0_ADD_7x7_fast_I32_Y_0 : AX1D
      port map(A => N165_1, B => N80, C => \un18_ready0_1[4]\, Y
         => \un18_ready0[4]\);
    
    un6_waddr_vect_s_I_16 : AND3
      port map(A => \data_mem_addr_w_0[0]\, B => 
        \data_mem_addr_w_0[1]\, C => \data_mem_addr_w_0[2]\, Y
         => \DWACT_FINC_E[0]\);
    
    un3_ready_0_0_0_ADD_5x5_fast_I18_Y_0 : XNOR2
      port map(A => N_6, B => N_89_i, Y => \un3_ready0[4]\);
    
    un18_ready_1_16_ADD_5x5_fast_I11_un1_Y : OR3C
      port map(A => N81, B => N77, C => N98, Y => I11_un1_Y);
    
    \Waddr_vect_RNIVOFL[0]\ : OR3A
      port map(A => \data_mem_wen_i_0[0]\, B => N_164, C => 
        \data_mem_addr_w_0[0]\, Y => N_157);
    
    sFull_RNO_1 : XA1
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \un8_waddr_vect_s[1]\, C => sFull_RNO_5_3, Y => 
        un5_sfull_s_4_1);
    
    \ready_gen.un12_ready_0_I_3\ : NOR2A
      port map(A => \data_mem_addr_r_0[0]\, B => 
        \data_mem_addr_w_0[0]\, Y => N_6_0);
    
    \Waddr_vect_RNIB0LI2[1]\ : NOR3C
      port map(A => N_149, B => data_addr_w_iv_i_2(1), C => N_150, 
        Y => data_addr_w_iv_i_4(1));
    
    un18_ready_1_16_ADD_5x5_fast_I0_CO1 : XA1B
      port map(A => \data_mem_addr_r_0[2]\, B => 
        \data_mem_addr_w_0[2]\, C => N_84_1, Y => N77);
    
    \Raddr_vect[3]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[0]\, Q => 
        \data_mem_addr_r_0[3]\);
    
    sFull_RNO_4 : OR2B
      port map(A => I_5_13, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[1]\);
    
    \Raddr_vect_RNI7G73_0[4]\ : NOR2A
      port map(A => \data_mem_addr_r_0[4]\, B => 
        \data_mem_addr_w_0[4]\, Y => N_75);
    
    sEmpty_RNO_5 : XNOR2
      port map(A => \un10_raddr_vect_s[2]\, B => 
        \data_mem_addr_w_0[2]\, Y => sEmpty_RNO_5_1);
    
    \Raddr_vect_RNI9B352[3]\ : OR2A
      port map(A => \data_mem_ren_i_0[0]\, B => 
        \data_mem_addr_r_0[3]\, Y => N_49);
    
    un3_ready_0_0_0_ADD_5x5_fast_I12_Y_i_a3 : AOI1
      port map(A => ADD_5x5_fast_I9_Y_i_o2_0, B => Waddr_vect_c1, 
        C => \data_mem_addr_r_0[2]\, Y => N_17);
    
    \Raddr_vect_RNI7G73[4]\ : XNOR2
      port map(A => \data_mem_addr_w_0[4]\, B => 
        \data_mem_addr_r_0[4]\, Y => N_89_i);
    
    \Raddr_vect_RNIM38B[4]\ : NOR2B
      port map(A => I_5_14, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[1]\);
    
    un8_raddr_vect_s_I_19 : NOR2B
      port map(A => \data_mem_addr_r_0[3]\, B => 
        \DWACT_FINC_E_0[0]\, Y => N_4_0);
    
    un3_ready_1_1_0_SUM2_0_0 : XOR2
      port map(A => N_89_i, B => N_109, Y => SUM2_0_0);
    
    \Raddr_vect[4]\ : DFN1E1C0
      port map(D => \un10_raddr_vect_s[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \data_mem_ren_i_0[0]\, Q => 
        \data_mem_addr_r_0[4]\);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_12, B => \data_mem_addr_w_0[2]\, Y => 
        I_9_13);
    
    \ready_gen.un12_ready_0_I_5\ : AO1C
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \data_mem_addr_w_0[1]\, C => N_6_0, Y => N_8);
    
    \ready_gen.un12_ready_0_I_1\ : OR2A
      port map(A => \data_mem_addr_r_0[1]\, B => 
        \data_mem_addr_w_0[1]\, Y => N_4_1);
    
    sEmpty_RNO_1 : NOR2B
      port map(A => \sEmpty\, B => data_wen(0), Y => un1_sempty_s);
    
    \Raddr_vect_RNICK9Q4[2]\ : NOR3C
      port map(A => data_addr_r_iv_i_1(2), B => 
        data_addr_r_iv_i_0(2), C => N_57, Y => 
        data_addr_r_iv_i_3(2));
    
    \Waddr_vect_RNI9473[3]\ : NOR2
      port map(A => \data_mem_addr_w_0[3]\, B => 
        \data_mem_addr_w_0[2]\, Y => un1_waddr_vect_slto3_0);
    
    un8_raddr_vect_s_I_20 : XOR2
      port map(A => N_4_0, B => \data_mem_addr_r_0[4]\, Y => 
        I_20_6);
    
    \ready_gen.un12_ready_0_I_4\ : OR2A
      port map(A => \data_mem_addr_r_0[4]\, B => 
        \data_mem_addr_w_0[4]\, Y => N_7);
    
    \Raddr_vect_RNI709Q4[1]\ : NOR3C
      port map(A => data_addr_r_iv_i_1(1), B => 
        data_addr_r_iv_i_0(1), C => N_65, Y => 
        data_addr_r_iv_i_3(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ4 is

    port( time_mem_ren_i_0_1   : in    std_logic;
          time_wen             : in    std_logic_vector(0 to 0);
          time_ren             : in    std_logic_vector(0 to 0);
          data_addr_w_0_iv_i_1 : out   std_logic_vector(5 to 5);
          Waddr_vect_RNILN58   : in    std_logic_vector(0 to 0);
          Waddr_vect_RNINV58   : in    std_logic_vector(2 to 2);
          Waddr_vect_RNI64MA   : in    std_logic_vector(2 to 2);
          data_addr_w_iv_i_2_0 : out   std_logic;
          data_addr_w_iv_i_2_2 : out   std_logic;
          time_mem_wen_i_0     : out   std_logic_vector(0 to 0);
          data_addr_r_0_iv_i_1 : in    std_logic_vector(5 to 5);
          data_addr_r_0_iv_i_2 : out   std_logic_vector(5 to 5);
          Raddr_vect_RNI8J9L   : in    std_logic_vector(2 to 2);
          data_addr_r_iv_i_0   : out   std_logic_vector(4 downto 0);
          data_addr_w_iv_i_1_0 : out   std_logic;
          data_addr_w_iv_i_1_3 : out   std_logic;
          data_addr_w_iv_i_1_1 : out   std_logic;
          HRESETn_c            : in    std_logic;
          HCLK_c               : in    std_logic;
          N_77                 : out   std_logic;
          sFull_RNI9VRD        : in    std_logic;
          N_140                : in    std_logic;
          sFull_RNIPQBB_0      : in    std_logic;
          N_122                : in    std_logic;
          N_124                : in    std_logic;
          sFull_RNI9VRD_0      : in    std_logic;
          N_146                : in    std_logic;
          N_70                 : in    std_logic;
          sEmpty_RNI5EFO_0     : in    std_logic;
          N_33                 : in    std_logic;
          N_62                 : in    std_logic;
          N_155                : in    std_logic;
          sFull_RNI9VRD_1      : in    std_logic;
          N_147                : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ4;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ4 is 

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \time_mem_addr_r_0[4]\, \Raddr_vect[2]_net_1\, 
        \Raddr_vect[3]_net_1\, N_4, \time_mem_addr_w_0[4]\, 
        \Waddr_vect[2]_net_1\, \Waddr_vect[3]_net_1\, N_4_0, N_7, 
        \time_mem_addr_r_0[1]\, \time_mem_addr_r_0[0]\, N_7_0, 
        \time_mem_addr_w_0[1]\, \time_mem_addr_w_0[0]\, 
        \data_addr_w_iv_i_0[1]\, \data_addr_w_iv_i_0[3]\, 
        \data_addr_w_iv_i_0[0]\, \time_mem_ren_i_0[0]\, 
        \time_mem_addr_r_0[3]\, \sEmpty_RNI2EFO\, 
        \data_addr_w_iv_i_0[4]\, \time_mem_wen_i_0[0]\, 
        \time_mem_addr_w_0[3]\, \data_addr_w_iv_i_0[2]\, 
        \sFull_RNIBMR8\, un7_sempty_s_3, \sEmpty_RNO_3\, 
        \sEmpty_RNO_4\, un7_sempty_s_0, un7_sempty_s_2, 
        \un10_raddr_vect_s[3]\, \un10_raddr_vect_s[0]\, 
        un5_sfull_s_2, \un8_waddr_vect_s[3]\, un5_sfull_s_1, 
        \un8_waddr_vect_s[1]\, \sFull_RNO_5\, un5_sfull_s_0, 
        \un8_waddr_vect_s[0]\, un2_raddr_vect_slt3, 
        un1_waddr_vect_slt3, un5_sfull_s, Raddr_vect_n3, 
        Raddr_vect_7_0, Waddr_vect_n3, Waddr_vect_15_0, 
        Raddr_vect_n2, un2_raddr_vect_s, Raddr_vect_n2_tz, 
        Waddr_vect_n2, un1_waddr_vect_s, Waddr_vect_n2_tz, 
        \sEmpty\, un2_sempty_s, \sFull\, \sEmpty_RNO_0\, 
        \sFull_RNO_0\, I_13_6, I_5_5, I_13_5, I_5_6, I_9_6, I_9_5, 
        Raddr_vect_n1_i, Raddr_vect_e2, Raddr_vect_e1, 
        Raddr_vect_e0, Waddr_vect_n1_i, Waddr_vect_e2, 
        Waddr_vect_e1, Waddr_vect_e0, N_4_1, N_4_2, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 

    time_mem_wen_i_0(0) <= \time_mem_wen_i_0[0]\;

    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_w_0[1]\, B => 
        \time_mem_addr_w_0[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_addr_w_0[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        N_4_1);
    
    sFull_RNI8KFI1 : NOR3C
      port map(A => sFull_RNI9VRD_0, B => \data_addr_w_iv_i_0[4]\, 
        C => N_124, Y => data_addr_w_iv_i_2_2);
    
    \Waddr_vect_RNI4JHO[1]\ : AND2
      port map(A => N_147, B => \data_addr_w_iv_i_0[1]\, Y => 
        data_addr_w_iv_i_1_1);
    
    \Raddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_r_0[1]\, B => 
        \time_mem_addr_r_0[0]\, C => un2_raddr_vect_s, Y => 
        Raddr_vect_n1_i);
    
    sEmpty_RNI2EFO : OR2
      port map(A => \time_mem_ren_i_0[0]\, B => N_4, Y => 
        \sEmpty_RNI2EFO\);
    
    \Waddr_vect_RNITOG9[1]\ : OR3
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_addr_w_0[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        un1_waddr_vect_slt3);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_w_0[1]\, B => 
        \time_mem_addr_w_0[0]\, Y => N_7_0);
    
    sEmpty_RNO : AO1
      port map(A => un7_sempty_s_3, B => un7_sempty_s_2, C => 
        un2_sempty_s, Y => \sEmpty_RNO_0\);
    
    \Raddr_vect[1]\ : DFN1C0
      port map(D => Raddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_0[1]\);
    
    \Waddr_vect[3]\ : DFN1E0C0
      port map(D => Waddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_wen_i_0[0]\, Q => 
        \Waddr_vect[3]_net_1\);
    
    sFull_RNIBMR8 : OR2
      port map(A => \time_mem_wen_i_0[0]\, B => N_4_0, Y => 
        \sFull_RNIBMR8\);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_7, B => \Raddr_vect[2]_net_1\, Y => I_9_6);
    
    \Raddr_vect_RNICUIA1[1]\ : OA1
      port map(A => \time_mem_addr_r_0[1]\, B => 
        \time_mem_ren_i_0[0]\, C => N_62, Y => 
        data_addr_r_iv_i_0(1));
    
    sEmpty : DFN1P0
      port map(D => \sEmpty_RNO_0\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \sEmpty\);
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => \time_mem_wen_i_0[0]\, 
        C => \time_mem_addr_w_0[0]\, Y => Waddr_vect_e0);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Waddr_vect[2]_net_1\);
    
    sFull_RNIA4G2 : OR2
      port map(A => time_wen(0), B => \sFull\, Y => 
        \time_mem_wen_i_0[0]\);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \time_mem_addr_w_0[1]\, 
        S => \time_mem_wen_i_0[0]\, Y => Waddr_vect_e1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Waddr_vect_RNO_0[2]\ : OR2B
      port map(A => un1_waddr_vect_s, B => Waddr_vect_n2_tz, Y
         => Waddr_vect_n2);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_addr_w_0[1]\, Y => I_5_5);
    
    \Raddr_vect_RNO_0[2]\ : OR2B
      port map(A => un2_raddr_vect_s, B => Raddr_vect_n2_tz, Y
         => Raddr_vect_n2);
    
    sEmpty_RNINO741 : NOR2B
      port map(A => time_mem_ren_i_0_1, B => 
        \time_mem_ren_i_0[0]\, Y => N_77);
    
    \Waddr_vect_RNIVIRD[1]\ : OA1
      port map(A => \time_mem_addr_w_0[1]\, B => 
        \time_mem_wen_i_0[0]\, C => N_146, Y => 
        \data_addr_w_iv_i_0[1]\);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => Raddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_ren_i_0[0]\, Q => 
        \Raddr_vect[3]_net_1\);
    
    sEmpty_RNO_2 : NOR2B
      port map(A => time_wen(0), B => \sEmpty\, Y => un2_sempty_s);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_4_1, B => \Waddr_vect[3]_net_1\, Y => 
        I_13_5);
    
    sFull_RNO : AO1
      port map(A => time_ren(0), B => \sFull\, C => un5_sfull_s, 
        Y => \sFull_RNO_0\);
    
    sEmpty_RNIBS3I : OR2
      port map(A => time_ren(0), B => \sEmpty\, Y => 
        \time_mem_ren_i_0[0]\);
    
    \Raddr_vect_RNO[0]\ : AXOI7
      port map(A => un2_raddr_vect_s, B => \time_mem_ren_i_0[0]\, 
        C => \time_mem_addr_r_0[0]\, Y => Raddr_vect_e0);
    
    \Raddr_vect_RNO[1]\ : MX2A
      port map(A => Raddr_vect_n1_i, B => \time_mem_addr_r_0[1]\, 
        S => \time_mem_ren_i_0[0]\, Y => Raddr_vect_e1);
    
    \Raddr_vect_RNIAMIA1[0]\ : OA1
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_ren_i_0[0]\, C => N_70, Y => 
        data_addr_r_iv_i_0(0));
    
    sFull_RNO_4 : OR2B
      port map(A => I_5_5, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[1]\);
    
    sFull_RNO_6 : OR2A
      port map(A => un1_waddr_vect_s, B => \time_mem_addr_w_0[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    sEmpty_RNO_3 : AX1E
      port map(A => un2_raddr_vect_s, B => I_9_6, C => 
        \Waddr_vect[2]_net_1\, Y => \sEmpty_RNO_3\);
    
    sEmpty_RNI7SUG1_0 : OA1
      port map(A => \time_mem_addr_r_0[3]\, B => 
        \time_mem_ren_i_0[0]\, C => sEmpty_RNI5EFO_0, Y => 
        data_addr_r_iv_i_0(3));
    
    \Raddr_vect[2]\ : DFN1C0
      port map(D => Raddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Raddr_vect[2]_net_1\);
    
    \Raddr_vect_RNIE6JA1[2]\ : OA1A
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \time_mem_ren_i_0[0]\, C => Raddr_vect_RNI8J9L(2), Y => 
        data_addr_r_iv_i_0(2));
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_0[0]\);
    
    sFull_RNO_5 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_5, C => 
        \Raddr_vect[2]_net_1\, Y => \sFull_RNO_5\);
    
    sFull_RNI4H7K : OA1B
      port map(A => \time_mem_addr_w_0[4]\, B => 
        \time_mem_wen_i_0[0]\, C => N_122, Y => 
        \data_addr_w_iv_i_0[4]\);
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => \Waddr_vect[2]_net_1\, S
         => \time_mem_wen_i_0[0]\, Y => Waddr_vect_e2);
    
    sEmpty_RNO_4 : AX1E
      port map(A => un2_raddr_vect_s, B => I_5_6, C => 
        \time_mem_addr_w_0[1]\, Y => \sEmpty_RNO_4\);
    
    sFull_RNO_3 : XA1
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \un8_waddr_vect_s[3]\, C => time_ren(0), Y => 
        un5_sfull_s_2);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => \sEmpty_RNO_3\, B => \sEmpty_RNO_4\, C => 
        un7_sempty_s_0, Y => un7_sempty_s_3);
    
    \Waddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_addr_w_0[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_n2_tz);
    
    un25_mem_addr_ren_I_8 : OR2B
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_0[4]\);
    
    sFull_RNIDG321 : NOR3B
      port map(A => \sFull_RNIBMR8\, B => sFull_RNI9VRD, C => 
        N_122, Y => data_addr_w_0_iv_i_1(5));
    
    \Waddr_vect_RNI1RRD[2]\ : OA1A
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \time_mem_wen_i_0[0]\, C => Waddr_vect_RNINV58(2), Y => 
        \data_addr_w_iv_i_0[2]\);
    
    \Raddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_addr_r_0[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        Raddr_vect_n2_tz);
    
    un25_mem_addr_ren_I_12 : NOR2B
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \Raddr_vect[2]_net_1\, Y => N_4);
    
    sEmpty_RNO_7 : OR2A
      port map(A => un2_raddr_vect_s, B => \time_mem_addr_r_0[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Raddr_vect_RNO[2]\ : MX2A
      port map(A => Raddr_vect_n2, B => \Raddr_vect[2]_net_1\, S
         => \time_mem_ren_i_0[0]\, Y => Raddr_vect_e2);
    
    \Raddr_vect[0]\ : DFN1C0
      port map(D => Raddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_0[0]\);
    
    sEmpty_RNI7SUG1 : OA1B
      port map(A => \time_mem_addr_r_0[4]\, B => 
        \time_mem_ren_i_0[0]\, C => N_33, Y => 
        data_addr_r_iv_i_0(4));
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_r_0[1]\, B => 
        \time_mem_addr_r_0[0]\, Y => N_7);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_7_0, B => \Waddr_vect[2]_net_1\, Y => I_9_5);
    
    \Waddr_vect_RNIU7O51[2]\ : NOR3C
      port map(A => Waddr_vect_RNI64MA(2), B => 
        \data_addr_w_iv_i_0[2]\, C => N_140, Y => 
        data_addr_w_iv_i_2_0);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_4_2, B => \Raddr_vect[3]_net_1\, Y => 
        I_13_6);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_addr_r_0[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        N_4_2);
    
    sFull_RNIDG321_0 : AND2
      port map(A => sFull_RNI9VRD_1, B => \data_addr_w_iv_i_0[3]\, 
        Y => data_addr_w_iv_i_1_3);
    
    sEmpty_RNO_1 : XA1B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \un10_raddr_vect_s[3]\, C => time_ren(0), Y => 
        un7_sempty_s_2);
    
    sFull_RNO_1 : XA1
      port map(A => \un8_waddr_vect_s[1]\, B => 
        \time_mem_addr_r_0[1]\, C => \sFull_RNO_5\, Y => 
        un5_sfull_s_1);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_addr_r_0[1]\, Y => I_5_6);
    
    \Raddr_vect_RNIEOG9[1]\ : OR3
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_addr_r_0[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        un2_raddr_vect_slt3);
    
    \Waddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_addr_w_0[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_15_0);
    
    sFull_RNO_7 : OR2B
      port map(A => I_13_5, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    \Waddr_vect_RNIUJMC[3]\ : OR2B
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, Y => un1_waddr_vect_s);
    
    \Raddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_r_0[0]\, B => 
        \time_mem_addr_r_0[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        Raddr_vect_7_0);
    
    sEmpty_RNIQOT13 : NOR3B
      port map(A => \sEmpty_RNI2EFO\, B => 
        data_addr_r_0_iv_i_1(5), C => N_33, Y => 
        data_addr_r_0_iv_i_2(5));
    
    un29_mem_addr_wen_I_8 : OR2B
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_0[4]\);
    
    un25_mem_addr_ren_I_5 : XOR2
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_0[3]\);
    
    \Waddr_vect_RNO[3]\ : AXOI1
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, C => Waddr_vect_15_0, Y => 
        Waddr_vect_n3);
    
    sFull_RNO_0 : NOR3C
      port map(A => un5_sfull_s_1, B => un5_sfull_s_0, C => 
        un5_sfull_s_2, Y => un5_sfull_s);
    
    sEmpty_RNO_6 : OR2B
      port map(A => I_13_6, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    un29_mem_addr_wen_I_5 : XOR2
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_0[3]\);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO_0\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \Waddr_vect_RNITARD[0]\ : OA1
      port map(A => \time_mem_addr_w_0[0]\, B => 
        \time_mem_wen_i_0[0]\, C => Waddr_vect_RNILN58(0), Y => 
        \data_addr_w_iv_i_0[0]\);
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_0[1]\);
    
    un29_mem_addr_wen_I_12 : NOR2B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \Waddr_vect[2]_net_1\, Y => N_4_0);
    
    sFull_RNO_2 : XA1B
      port map(A => \un8_waddr_vect_s[0]\, B => 
        \time_mem_addr_r_0[0]\, C => time_wen(0), Y => 
        un5_sfull_s_0);
    
    sFull_RNI4H7K_0 : OA1
      port map(A => \time_mem_addr_w_0[3]\, B => 
        \time_mem_wen_i_0[0]\, C => sFull_RNIPQBB_0, Y => 
        \data_addr_w_iv_i_0[3]\);
    
    sEmpty_RNO_5 : XA1
      port map(A => \un10_raddr_vect_s[0]\, B => 
        \time_mem_addr_w_0[0]\, C => time_wen(0), Y => 
        un7_sempty_s_0);
    
    \Raddr_vect_RNO[3]\ : AXOI1
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, C => Raddr_vect_7_0, Y => 
        Raddr_vect_n3);
    
    \Raddr_vect_RNIAJMC[3]\ : OR2B
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, Y => un2_raddr_vect_s);
    
    \Waddr_vect_RNI17HO[0]\ : AND2
      port map(A => N_155, B => \data_addr_w_iv_i_0[0]\, Y => 
        data_addr_w_iv_i_1_0);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_ctrlZ6 is

    port( Waddr_vect_RNI64MA       : out   std_logic_vector(2 to 2);
          data_addr_w_1_iv_i_s_0_0 : in    std_logic_vector(6 to 6);
          time_wen                 : in    std_logic_vector(2 to 2);
          data_addr_r_0_iv_i_1     : out   std_logic_vector(5 to 5);
          data_addr_r_1_iv_i_s_1   : out   std_logic_vector(6 to 6);
          time_mem_ren_i_0_1       : in    std_logic;
          data_addr_r_iv_i_a2_0    : out   std_logic_vector(4 to 4);
          data_addr_r_iv_i_1       : out   std_logic_vector(4 downto 0);
          time_ren                 : in    std_logic_vector(2 to 2);
          time_ren_1z              : in    std_logic;
          HRESETn_c                : in    std_logic;
          HCLK_c                   : in    std_logic;
          sFull_RNI9VRD_0          : out   std_logic;
          N_147                    : out   std_logic;
          sFull_RNI9VRD_1          : out   std_logic;
          sFull_RNI9VRD            : out   std_logic;
          un13_time_write          : in    std_logic;
          N_163                    : out   std_logic;
          N_155                    : out   std_logic;
          N_162                    : in    std_logic;
          sFull_RNIU5GK1           : out   std_logic;
          N_29                     : in    std_logic;
          N_30_1                   : in    std_logic;
          N_72                     : in    std_logic;
          N_56                     : in    std_logic;
          N_48                     : in    std_logic;
          N_35                     : in    std_logic;
          N_64                     : in    std_logic
        );

end lpp_waveform_fifo_ctrlZ6;

architecture DEF_ARCH of lpp_waveform_fifo_ctrlZ6 is 

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \time_mem_addr_r_2[4]\, \Raddr_vect[2]_net_1\, 
        \Raddr_vect[3]_net_1\, N_4, \time_mem_addr_w_2[4]\, 
        \Waddr_vect[2]_net_1\, \Waddr_vect[3]_net_1\, N_4_0, N_7, 
        \time_mem_addr_r_2[1]\, \time_mem_addr_r_2[0]\, N_7_0, 
        \time_mem_addr_w_2[1]\, \time_mem_addr_w_2[0]\, 
        \un2_sfull_s_3_0\, \un8_waddr_vect_s[3]\, 
        \un10_sempty_s_3_0\, \un10_raddr_vect_s[3]\, 
        un5_sfull_s_2, un7_sempty_s_2, \time_mem_ren_i_0[2]\, 
        \time_mem_addr_r_2[3]\, un5_sfull_s_3, \sFull_RNO_3\, 
        \sFull_RNO_4\, un5_sfull_s_0, \un8_waddr_vect_s[0]\, 
        un7_sempty_s_3, sEmpty_RNO_3_0, sEmpty_RNO_4_0, 
        un7_sempty_s_0, \un10_raddr_vect_s[0]\, 
        un2_raddr_vect_slt3, \time_mem_wen_i_0[2]\, 
        un1_waddr_vect_slt3, Raddr_vect_n3, Raddr_vect_7_0, 
        Waddr_vect_n3, Waddr_vect_15_0, Raddr_vect_c1, 
        Raddr_vect_n2, un2_raddr_vect_s, Waddr_vect_n2, 
        un1_waddr_vect_s, Waddr_vect_n2_tz, I_13_7, I_9_7, I_5_7, 
        I_9_8, I_5_8, Raddr_vect_n1_i, N_50, Raddr_vect_e2, 
        Raddr_vect_e1, Raddr_vect_e0, I_13_8, \sFull_RNO_1\, 
        un8_sfull_s, \sEmpty_RNO_1\, un2_sempty_s, \sFull\, 
        \sEmpty\, Waddr_vect_n1_i, Waddr_vect_e2, Waddr_vect_e1, 
        Waddr_vect_e0, \time_mem_addr_w_2[3]\, N_4_1, N_4_2, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Waddr_vect_RNO_0[1]\ : XAI1
      port map(A => \time_mem_addr_w_2[1]\, B => 
        \time_mem_addr_w_2[0]\, C => un1_waddr_vect_s, Y => 
        Waddr_vect_n1_i);
    
    un6_waddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_w_2[0]\, B => 
        \time_mem_addr_w_2[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        N_4_1);
    
    un37_mem_addr_ren_I_8 : OR2B
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_2[4]\);
    
    sEmpty_RNITO232 : NOR3C
      port map(A => N_30_1, B => \time_mem_ren_i_0[2]\, C => N_29, 
        Y => data_addr_r_1_iv_i_s_1(6));
    
    \Raddr_vect_RNO_0[1]\ : AX1C
      port map(A => un2_raddr_vect_s, B => \time_mem_addr_r_2[1]\, 
        C => N_50, Y => Raddr_vect_n1_i);
    
    \Waddr_vect_RNI4SLA[0]\ : OR3
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => 
        \time_mem_addr_w_2[0]\, Y => N_155);
    
    \sFull_RNI9VRD_1\ : OR3
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => 
        \time_mem_addr_w_2[3]\, Y => sFull_RNI9VRD_1);
    
    \sFull_RNI9VRD_0\ : OR3
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => 
        \time_mem_addr_w_2[4]\, Y => sFull_RNI9VRD_0);
    
    un6_waddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_w_2[1]\, B => 
        \time_mem_addr_w_2[0]\, Y => N_7_0);
    
    sEmpty_RNO : AO1
      port map(A => un7_sempty_s_3, B => un7_sempty_s_2, C => 
        un2_sempty_s, Y => \sEmpty_RNO_1\);
    
    \Raddr_vect[1]\ : DFN1C0
      port map(D => Raddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_2[1]\);
    
    \Waddr_vect[3]\ : DFN1E0C0
      port map(D => Waddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_wen_i_0[2]\, Q => 
        \Waddr_vect[3]_net_1\);
    
    \Raddr_vect_RNIKOG9[1]\ : OR3
      port map(A => \time_mem_addr_r_2[0]\, B => 
        \time_mem_addr_r_2[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        un2_raddr_vect_slt3);
    
    un8_raddr_vect_s_I_9 : XOR2
      port map(A => N_7, B => \Raddr_vect[2]_net_1\, Y => I_9_8);
    
    un2_sfull_s_3_0_RNO : OR2B
      port map(A => I_13_7, B => un1_waddr_vect_s, Y => 
        \un8_waddr_vect_s[3]\);
    
    sEmpty : DFN1P0
      port map(D => \sEmpty_RNO_1\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \sEmpty\);
    
    \Waddr_vect_RNO[0]\ : AXOI7
      port map(A => un1_waddr_vect_s, B => \time_mem_wen_i_0[2]\, 
        C => \time_mem_addr_w_2[0]\, Y => Waddr_vect_e0);
    
    \Waddr_vect[2]\ : DFN1C0
      port map(D => Waddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Waddr_vect[2]_net_1\);
    
    \Waddr_vect_RNO[1]\ : MX2A
      port map(A => Waddr_vect_n1_i, B => \time_mem_addr_w_2[1]\, 
        S => \time_mem_wen_i_0[2]\, Y => Waddr_vect_e1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Waddr_vect_RNO_0[2]\ : OR2B
      port map(A => un1_waddr_vect_s, B => Waddr_vect_n2_tz, Y
         => Waddr_vect_n2);
    
    un6_waddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_w_2[0]\, B => 
        \time_mem_addr_w_2[1]\, Y => I_5_7);
    
    \sFull_RNI9VRD\ : OR3
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => N_4_0, 
        Y => sFull_RNI9VRD);
    
    \Raddr_vect_RNO_0[2]\ : XAI1
      port map(A => \Raddr_vect[2]_net_1\, B => Raddr_vect_c1, C
         => un2_raddr_vect_s, Y => Raddr_vect_n2);
    
    \Raddr_vect[3]\ : DFN1E0C0
      port map(D => Raddr_vect_n3, CLK => HCLK_c, CLR => 
        HRESETn_c, E => \time_mem_ren_i_0[2]\, Q => 
        \Raddr_vect[3]_net_1\);
    
    \Waddr_vect_RNI64MA[2]\ : OR3A
      port map(A => \Waddr_vect[2]_net_1\, B => N_162, C => 
        \time_mem_wen_i_0[2]\, Y => Waddr_vect_RNI64MA(2));
    
    sEmpty_RNO_2 : NOR2B
      port map(A => time_wen(2), B => \sEmpty\, Y => un2_sempty_s);
    
    un6_waddr_vect_s_I_13 : XOR2
      port map(A => N_4_1, B => \Waddr_vect[3]_net_1\, Y => 
        I_13_7);
    
    un2_sfull_s_3_0 : XOR2
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \un8_waddr_vect_s[3]\, Y => \un2_sfull_s_3_0\);
    
    sFull_RNO : AO1
      port map(A => un5_sfull_s_3, B => un5_sfull_s_2, C => 
        un8_sfull_s, Y => \sFull_RNO_1\);
    
    \Raddr_vect_RNO[0]\ : AXOI7
      port map(A => un2_raddr_vect_s, B => \time_mem_ren_i_0[2]\, 
        C => \time_mem_addr_r_2[0]\, Y => Raddr_vect_e0);
    
    \Raddr_vect_RNO[1]\ : MX2A
      port map(A => Raddr_vect_n1_i, B => \time_mem_addr_r_2[1]\, 
        S => \time_mem_ren_i_0[2]\, Y => Raddr_vect_e1);
    
    sFull_RNO_4 : AX1E
      port map(A => un1_waddr_vect_s, B => I_5_7, C => 
        \time_mem_addr_r_2[1]\, Y => \sFull_RNO_4\);
    
    sFull_RNO_6 : OR2A
      port map(A => un1_waddr_vect_s, B => \time_mem_addr_w_2[0]\, 
        Y => \un8_waddr_vect_s[0]\);
    
    sEmpty_RNO_3 : AX1E
      port map(A => un2_raddr_vect_s, B => I_9_8, C => 
        \Waddr_vect[2]_net_1\, Y => sEmpty_RNO_3_0);
    
    \Raddr_vect[2]\ : DFN1C0
      port map(D => Raddr_vect_e2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \Raddr_vect[2]_net_1\);
    
    sEmpty_RNIJSUG1_0 : OA1
      port map(A => N_4, B => \time_mem_ren_i_0[2]\, C => N_35, Y
         => data_addr_r_0_iv_i_1(5));
    
    \Waddr_vect[0]\ : DFN1C0
      port map(D => Waddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_2[0]\);
    
    sFull_RNO_5 : XA1B
      port map(A => \un8_waddr_vect_s[0]\, B => 
        \time_mem_addr_r_2[0]\, C => time_wen(2), Y => 
        un5_sfull_s_0);
    
    \Waddr_vect_RNO[2]\ : MX2A
      port map(A => Waddr_vect_n2, B => \Waddr_vect[2]_net_1\, S
         => \time_mem_wen_i_0[2]\, Y => Waddr_vect_e2);
    
    sEmpty_RNO_4 : AX1E
      port map(A => un2_raddr_vect_s, B => I_5_8, C => 
        \time_mem_addr_w_2[1]\, Y => sEmpty_RNO_4_0);
    
    \Raddr_vect_RNIN1B6[1]\ : NOR2B
      port map(A => \time_mem_addr_r_2[1]\, B => 
        \time_mem_addr_r_2[0]\, Y => Raddr_vect_c1);
    
    \Waddr_vect_RNI3PG9[1]\ : OR3
      port map(A => \time_mem_addr_w_2[0]\, B => 
        \time_mem_addr_w_2[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        un1_waddr_vect_slt3);
    
    un10_sempty_s_3_0 : XOR2
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \un10_raddr_vect_s[3]\, Y => \un10_sempty_s_3_0\);
    
    \Raddr_vect_RNIIMIA1[0]\ : OA1
      port map(A => \time_mem_addr_r_2[0]\, B => 
        \time_mem_ren_i_0[2]\, C => N_72, Y => 
        data_addr_r_iv_i_1(0));
    
    un43_mem_addr_wen_I_12 : NOR2B
      port map(A => \Waddr_vect[3]_net_1\, B => 
        \Waddr_vect[2]_net_1\, Y => N_4_0);
    
    sFull_RNO_3 : AX1E
      port map(A => un1_waddr_vect_s, B => I_9_7, C => 
        \Raddr_vect[2]_net_1\, Y => \sFull_RNO_3\);
    
    sEmpty_RNO_0 : NOR3C
      port map(A => sEmpty_RNO_3_0, B => sEmpty_RNO_4_0, C => 
        un7_sempty_s_0, Y => un7_sempty_s_3);
    
    \Waddr_vect_RNO_1[2]\ : AX1C
      port map(A => \time_mem_addr_w_2[0]\, B => 
        \time_mem_addr_w_2[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_n2_tz);
    
    un43_mem_addr_wen_I_8 : OR2B
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_2[4]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Raddr_vect_RNO[2]\ : MX2A
      port map(A => Raddr_vect_n2, B => \Raddr_vect[2]_net_1\, S
         => \time_mem_ren_i_0[2]\, Y => Raddr_vect_e2);
    
    \Raddr_vect[0]\ : DFN1C0
      port map(D => Raddr_vect_e0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_r_2[0]\);
    
    \Waddr_vect_RNI50MA[1]\ : OR3
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => 
        \time_mem_addr_w_2[1]\, Y => N_147);
    
    sEmpty_RNIRO741 : NOR2B
      port map(A => time_mem_ren_i_0_1, B => 
        \time_mem_ren_i_0[2]\, Y => data_addr_r_iv_i_a2_0(4));
    
    un8_raddr_vect_s_I_8 : NOR2B
      port map(A => \time_mem_addr_r_2[1]\, B => 
        \time_mem_addr_r_2[0]\, Y => N_7);
    
    un10_sempty_s_3_0_RNO : OR2B
      port map(A => I_13_8, B => un2_raddr_vect_s, Y => 
        \un10_raddr_vect_s[3]\);
    
    un6_waddr_vect_s_I_9 : XOR2
      port map(A => N_7_0, B => \Waddr_vect[2]_net_1\, Y => I_9_7);
    
    un8_raddr_vect_s_I_13 : XOR2
      port map(A => N_4_2, B => \Raddr_vect[3]_net_1\, Y => 
        I_13_8);
    
    un8_raddr_vect_s_I_12 : AND3
      port map(A => \time_mem_addr_r_2[0]\, B => 
        \time_mem_addr_r_2[1]\, C => \Raddr_vect[2]_net_1\, Y => 
        N_4_2);
    
    \Raddr_vect_RNIKUIA1[1]\ : OA1
      port map(A => \time_mem_addr_r_2[1]\, B => 
        \time_mem_ren_i_0[2]\, C => N_64, Y => 
        data_addr_r_iv_i_1(1));
    
    sEmpty_RNO_1 : NOR2A
      port map(A => \un10_sempty_s_3_0\, B => time_ren(2), Y => 
        un7_sempty_s_2);
    
    \Raddr_vect_RNIM6JA1[2]\ : OA1A
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \time_mem_ren_i_0[2]\, C => N_56, Y => 
        data_addr_r_iv_i_1(2));
    
    sEmpty_RNIDS3I : OR3A
      port map(A => time_ren_1z, B => un13_time_write, C => 
        \sEmpty\, Y => \time_mem_ren_i_0[2]\);
    
    sFull_RNO_1 : AND2
      port map(A => time_ren(2), B => \un2_sfull_s_3_0\, Y => 
        un5_sfull_s_2);
    
    un8_raddr_vect_s_I_5 : XOR2
      port map(A => \time_mem_addr_r_2[0]\, B => 
        \time_mem_addr_r_2[1]\, Y => I_5_8);
    
    un43_mem_addr_wen_I_5 : XOR2
      port map(A => \Waddr_vect[2]_net_1\, B => 
        \Waddr_vect[3]_net_1\, Y => \time_mem_addr_w_2[3]\);
    
    \Waddr_vect_RNI6KMC[3]\ : OR2B
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, Y => un1_waddr_vect_s);
    
    un37_mem_addr_ren_I_12 : NOR2B
      port map(A => \Raddr_vect[3]_net_1\, B => 
        \Raddr_vect[2]_net_1\, Y => N_4);
    
    \Waddr_vect_RNO_0[3]\ : OR3C
      port map(A => \time_mem_addr_w_2[0]\, B => 
        \time_mem_addr_w_2[1]\, C => \Waddr_vect[2]_net_1\, Y => 
        Waddr_vect_15_0);
    
    \Raddr_vect_RNO_0[3]\ : OR2B
      port map(A => Raddr_vect_c1, B => \Raddr_vect[2]_net_1\, Y
         => Raddr_vect_7_0);
    
    \Raddr_vect_RNIIJMC[3]\ : OR2B
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, Y => un2_raddr_vect_s);
    
    \Waddr_vect_RNO[3]\ : AXOI1
      port map(A => un1_waddr_vect_slt3, B => 
        \Waddr_vect[3]_net_1\, C => Waddr_vect_15_0, Y => 
        Waddr_vect_n3);
    
    sFull_RNI4DG7 : NOR2A
      port map(A => \time_mem_wen_i_0[2]\, B => N_162, Y => N_163);
    
    sFull_RNO_0 : NOR3C
      port map(A => \sFull_RNO_3\, B => \sFull_RNO_4\, C => 
        un5_sfull_s_0, Y => un5_sfull_s_3);
    
    sEmpty_RNO_6 : OR2A
      port map(A => un2_raddr_vect_s, B => \time_mem_addr_r_2[0]\, 
        Y => \un10_raddr_vect_s[0]\);
    
    un37_mem_addr_ren_I_5 : XOR2
      port map(A => \Raddr_vect[2]_net_1\, B => 
        \Raddr_vect[3]_net_1\, Y => \time_mem_addr_r_2[3]\);
    
    sEmpty_RNIJSUG1_1 : OA1
      port map(A => \time_mem_addr_r_2[4]\, B => 
        \time_mem_ren_i_0[2]\, C => N_35, Y => 
        data_addr_r_iv_i_1(4));
    
    \Raddr_vect_RNO_1[1]\ : OR2B
      port map(A => \time_mem_addr_r_2[0]\, B => un2_raddr_vect_s, 
        Y => N_50);
    
    sFull : DFN1C0
      port map(D => \sFull_RNO_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \sFull\);
    
    \sFull_RNIU5GK1\ : OAI1
      port map(A => N_162, B => \time_mem_wen_i_0[2]\, C => 
        data_addr_w_1_iv_i_s_0_0(6), Y => sFull_RNIU5GK1);
    
    sFull_RNIE4G2 : OR2
      port map(A => time_wen(2), B => \sFull\, Y => 
        \time_mem_wen_i_0[2]\);
    
    sEmpty_RNIJSUG1 : OA1
      port map(A => \time_mem_addr_r_2[3]\, B => 
        \time_mem_ren_i_0[2]\, C => N_48, Y => 
        data_addr_r_iv_i_1(3));
    
    \Waddr_vect[1]\ : DFN1C0
      port map(D => Waddr_vect_e1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \time_mem_addr_w_2[1]\);
    
    sFull_RNO_2 : OA1A
      port map(A => time_ren_1z, B => un13_time_write, C => 
        \sFull\, Y => un8_sfull_s);
    
    sEmpty_RNO_5 : XA1
      port map(A => \un10_raddr_vect_s[0]\, B => 
        \time_mem_addr_w_2[0]\, C => time_wen(2), Y => 
        un7_sempty_s_0);
    
    \Raddr_vect_RNO[3]\ : AXOI1
      port map(A => un2_raddr_vect_slt3, B => 
        \Raddr_vect[3]_net_1\, C => Raddr_vect_7_0, Y => 
        Raddr_vect_n3);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo is

    port( data_wen              : in    std_logic_vector(3 downto 0);
          data_ren              : in    std_logic_vector(3 downto 0);
          ready_i_0             : out   std_logic_vector(3 downto 0);
          time_ren              : in    std_logic_vector(3 downto 0);
          time_wen              : in    std_logic_vector(3 downto 0);
          wdata                 : in    std_logic_vector(31 downto 0);
          hwdata_c              : out   std_logic_vector(31 downto 0);
          time_ren_1z           : in    std_logic;
          data_ren_1z           : in    std_logic;
          un20_time_write       : in    std_logic;
          un13_time_write       : in    std_logic;
          HRESETn_c             : in    std_logic;
          lpp_waveform_fifo_VCC : in    std_logic;
          lpp_waveform_fifo_GND : in    std_logic;
          HCLK_c                : in    std_logic
        );

end lpp_waveform_fifo;

architecture DEF_ARCH of lpp_waveform_fifo is 

  component lpp_waveform_fifo_ctrlZ1
    port( ready_i_0             : out   std_logic_vector(1 to 1);
          Raddr_vect_RNICA1PH   : out   std_logic_vector(1 to 1);
          data_mem_wen_i_0      : inout   std_logic_vector(2 downto 1);
          Raddr_vect_RNIIMQ5I   : out   std_logic_vector(4 to 4);
          Raddr_vect_RNIE6Q5I   : out   std_logic_vector(3 to 3);
          Raddr_vect_RNIKA2PH   : out   std_logic_vector(2 to 2);
          data_addr_r_iv_i_3    : in    std_logic_vector(4 downto 0) := (others => 'U');
          Raddr_vect_RNI4A0PH   : out   std_logic_vector(0 to 0);
          data_addr_r_iv_i_a2_2 : in    std_logic_vector(4 to 4) := (others => 'U');
          data_wen              : in    std_logic_vector(1 to 1) := (others => 'U');
          data_mem_ren_i_0      : inout   std_logic_vector(1 downto 0);
          data_ren              : in    std_logic_vector(1 to 1) := (others => 'U');
          data_ren_1z           : in    std_logic := 'U';
          HRESETn_c             : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U';
          N_166                 : out   std_logic;
          N_126                 : out   std_logic;
          N_150                 : out   std_logic;
          N_134                 : out   std_logic;
          N_142                 : out   std_logic;
          N_165                 : in    std_logic := 'U';
          N_158                 : out   std_logic;
          un20_time_write       : in    std_logic := 'U';
          N_68                  : in    std_logic := 'U';
          N_164                 : in    std_logic := 'U';
          N_120_i               : out   std_logic;
          N_44                  : in    std_logic := 'U';
          N_52                  : in    std_logic := 'U';
          N_60                  : in    std_logic := 'U';
          N_76                  : in    std_logic := 'U';
          N_86                  : out   std_logic;
          N_75                  : in    std_logic := 'U';
          N_59                  : in    std_logic := 'U';
          N_51                  : in    std_logic := 'U';
          N_43                  : in    std_logic := 'U';
          N_67                  : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component lpp_waveform_fifo_ctrlZ7
    port( time_mem_addr_w_3_i_0_1     : out   std_logic;
          data_addr_w_1_iv_i_a2_1_1_0 : in    std_logic_vector(6 to 6) := (others => 'U');
          data_addr_w_1_iv_i_s_0_0    : out   std_logic_vector(6 to 6);
          time_wen                    : in    std_logic_vector(3 to 3) := (others => 'U');
          time_ren                    : in    std_logic_vector(3 to 3) := (others => 'U');
          data_mem_ren_i_0            : in    std_logic_vector(1 to 1) := (others => 'U');
          time_mem_ren_i_0            : out   std_logic_vector(3 to 3);
          data_addr_r_1_iv_i_a9_1_1   : out   std_logic_vector(6 to 6);
          time_mem_addr_w_3           : out   std_logic_vector(1 downto 0);
          HRESETn_c                   : in    std_logic := 'U';
          HCLK_c                      : in    std_logic := 'U';
          N_124                       : out   std_logic;
          N_64                        : out   std_logic;
          N_140                       : out   std_logic;
          N_30_1                      : out   std_logic;
          N_89                        : out   std_logic;
          N_163                       : in    std_logic := 'U';
          N_164                       : out   std_logic;
          N_72                        : out   std_logic;
          N_56                        : out   std_logic;
          N_48                        : out   std_logic;
          N_35                        : out   std_logic;
          N_113                       : in    std_logic := 'U';
          N_162                       : in    std_logic := 'U';
          N_77                        : in    std_logic := 'U'
        );
  end component;

  component syncram_2pZ1
    port( hwdata_c            : out   std_logic_vector(31 downto 0);
          Raddr_vect_RNI4A0PH : in    std_logic_vector(0 to 0) := (others => 'U');
          Raddr_vect_RNICA1PH : in    std_logic_vector(1 to 1) := (others => 'U');
          Raddr_vect_RNIKA2PH : in    std_logic_vector(2 to 2) := (others => 'U');
          Raddr_vect_RNIE6Q5I : in    std_logic_vector(3 to 3) := (others => 'U');
          Raddr_vect_RNIIMQ5I : in    std_logic_vector(4 to 4) := (others => 'U');
          Waddr_vect_RNION355 : in    std_logic_vector(0 to 0) := (others => 'U');
          Waddr_vect_RNI0O455 : in    std_logic_vector(1 to 1) := (others => 'U');
          Waddr_vect_RNI394D5 : in    std_logic_vector(2 to 2) := (others => 'U');
          Waddr_vect_RNIJTNE5 : in    std_logic_vector(3 to 3) := (others => 'U');
          Waddr_vect_RNILLSP5 : in    std_logic_vector(4 to 4) := (others => 'U');
          wdata               : in    std_logic_vector(31 downto 0) := (others => 'U');
          HCLK_c              : in    std_logic := 'U';
          N_1_i_1             : in    std_logic := 'U';
          sEmpty_RNIE7T87     : in    std_logic := 'U';
          sEmpty_RNILSD08     : in    std_logic := 'U';
          sFull_RNIHL443      : in    std_logic := 'U';
          sFull_RNIU5GK1      : in    std_logic := 'U';
          syncram_2pZ1_GND    : in    std_logic := 'U';
          syncram_2pZ1_VCC    : in    std_logic := 'U';
          N_1_i_1_i           : in    std_logic := 'U'
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component lpp_waveform_fifo_ctrlZ2
    port( ready_i_0             : out   std_logic_vector(2 to 2);
          data_mem_wen_i_0      : out   std_logic_vector(2 to 2);
          data_ren              : in    std_logic_vector(2 to 2) := (others => 'U');
          Waddr_vect_RNI0O455   : out   std_logic_vector(1 to 1);
          Waddr_vect_RNILLSP5   : out   std_logic_vector(4 to 4);
          Waddr_vect_RNIJTNE5   : out   std_logic_vector(3 to 3);
          Waddr_vect_RNI394D5   : out   std_logic_vector(2 to 2);
          data_mem_ren_i_0_0    : in    std_logic := 'U';
          data_addr_r_0_iv_i_2  : in    std_logic_vector(5 to 5) := (others => 'U');
          data_addr_w_iv_i_4    : in    std_logic_vector(4 downto 0) := (others => 'U');
          Waddr_vect_RNION355   : out   std_logic_vector(0 to 0);
          data_wen              : in    std_logic_vector(2 to 2) := (others => 'U');
          data_addr_r_iv_i_a2_0 : in    std_logic_vector(4 to 4) := (others => 'U');
          data_addr_r_iv_i_a2_2 : out   std_logic_vector(4 to 4);
          HRESETn_c             : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U';
          N_67                  : out   std_logic;
          N_166                 : in    std_logic := 'U';
          N_75                  : out   std_logic;
          N_59                  : out   std_logic;
          N_51                  : out   std_logic;
          N_43                  : out   std_logic;
          N_152                 : in    std_logic := 'U';
          N_128                 : in    std_logic := 'U';
          N_136                 : in    std_logic := 'U';
          N_144                 : in    std_logic := 'U';
          sEmpty_RNIE7T87       : out   std_logic;
          N_160                 : in    std_logic := 'U';
          N_77                  : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_fifo_ctrlZ5
    port( time_mem_wen_i_0_0 : in    std_logic := 'U';
          Waddr_vect_RNINV58 : out   std_logic_vector(2 to 2);
          Waddr_vect_RNILN58 : out   std_logic_vector(0 to 0);
          Raddr_vect_RNI8J9L : out   std_logic_vector(2 to 2);
          time_mem_ren_i_0   : out   std_logic_vector(1 to 1);
          time_wen           : in    std_logic_vector(1 to 1) := (others => 'U');
          time_ren           : in    std_logic_vector(1 to 1) := (others => 'U');
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          N_146              : out   std_logic;
          N_162              : out   std_logic;
          N_113              : out   std_logic;
          N_122              : out   std_logic;
          sFull_RNIPQBB_0    : out   std_logic;
          N_62               : out   std_logic;
          N_70               : out   std_logic;
          sEmpty_RNI5EFO_0   : out   std_logic;
          N_33               : out   std_logic;
          N_29               : out   std_logic
        );
  end component;

  component lpp_waveform_fifo_ctrlZ3
    port( ready_i_0          : out   std_logic_vector(3 to 3);
          data_mem_wen_i_0_0 : in    std_logic := 'U';
          data_ren           : in    std_logic_vector(3 to 3) := (others => 'U');
          data_wen           : in    std_logic_vector(3 to 3) := (others => 'U');
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          N_128              : out   std_logic;
          N_152              : out   std_logic;
          N_136              : out   std_logic;
          N_68               : out   std_logic;
          N_144              : out   std_logic;
          N_166              : in    std_logic := 'U';
          N_160              : out   std_logic;
          N_76               : out   std_logic;
          N_60               : out   std_logic;
          N_52               : out   std_logic;
          N_86               : in    std_logic := 'U';
          N_44               : out   std_logic;
          N_1_i_1            : out   std_logic;
          N_1_i_1_i          : out   std_logic
        );
  end component;

  component lpp_waveform_fifo_ctrlZ0
    port( ready_i_0                   : out   std_logic_vector(0 to 0);
          data_ren                    : in    std_logic_vector(0 to 0) := (others => 'U');
          data_addr_w_0_iv_i_1        : in    std_logic_vector(5 to 5) := (others => 'U');
          data_addr_r_1_iv_i_s_1      : in    std_logic_vector(6 to 6) := (others => 'U');
          data_addr_r_1_iv_i_a9_1_1   : in    std_logic_vector(6 to 6) := (others => 'U');
          data_mem_ren_i_0            : out   std_logic_vector(0 to 0);
          data_mem_wen_i_0_1          : in    std_logic := 'U';
          data_addr_w_1_iv_i_a2_1_1_0 : out   std_logic_vector(6 to 6);
          data_addr_w_iv_i_2          : in    std_logic_vector(4 downto 0) := (others => 'U');
          data_addr_w_iv_i_4          : out   std_logic_vector(4 downto 0);
          data_wen                    : in    std_logic_vector(0 to 0) := (others => 'U');
          data_addr_r_iv_i_0          : in    std_logic_vector(4 downto 0) := (others => 'U');
          data_addr_r_iv_i_1          : in    std_logic_vector(4 downto 0) := (others => 'U');
          data_addr_r_iv_i_3          : out   std_logic_vector(4 downto 0);
          HRESETn_c                   : in    std_logic := 'U';
          HCLK_c                      : in    std_logic := 'U';
          N_165                       : out   std_logic;
          N_120_i                     : in    std_logic := 'U';
          sFull_RNIHL443              : out   std_logic;
          sEmpty_RNILSD08             : out   std_logic;
          N_124                       : in    std_logic := 'U';
          N_164                       : in    std_logic := 'U';
          N_158                       : in    std_logic := 'U';
          N_142                       : in    std_logic := 'U';
          N_134                       : in    std_logic := 'U';
          N_126                       : in    std_logic := 'U';
          N_150                       : in    std_logic := 'U'
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component lpp_waveform_fifo_ctrlZ4
    port( time_mem_ren_i_0_1   : in    std_logic := 'U';
          time_wen             : in    std_logic_vector(0 to 0) := (others => 'U');
          time_ren             : in    std_logic_vector(0 to 0) := (others => 'U');
          data_addr_w_0_iv_i_1 : out   std_logic_vector(5 to 5);
          Waddr_vect_RNILN58   : in    std_logic_vector(0 to 0) := (others => 'U');
          Waddr_vect_RNINV58   : in    std_logic_vector(2 to 2) := (others => 'U');
          Waddr_vect_RNI64MA   : in    std_logic_vector(2 to 2) := (others => 'U');
          data_addr_w_iv_i_2_0 : out   std_logic;
          data_addr_w_iv_i_2_2 : out   std_logic;
          time_mem_wen_i_0     : out   std_logic_vector(0 to 0);
          data_addr_r_0_iv_i_1 : in    std_logic_vector(5 to 5) := (others => 'U');
          data_addr_r_0_iv_i_2 : out   std_logic_vector(5 to 5);
          Raddr_vect_RNI8J9L   : in    std_logic_vector(2 to 2) := (others => 'U');
          data_addr_r_iv_i_0   : out   std_logic_vector(4 downto 0);
          data_addr_w_iv_i_1_0 : out   std_logic;
          data_addr_w_iv_i_1_3 : out   std_logic;
          data_addr_w_iv_i_1_1 : out   std_logic;
          HRESETn_c            : in    std_logic := 'U';
          HCLK_c               : in    std_logic := 'U';
          N_77                 : out   std_logic;
          sFull_RNI9VRD        : in    std_logic := 'U';
          N_140                : in    std_logic := 'U';
          sFull_RNIPQBB_0      : in    std_logic := 'U';
          N_122                : in    std_logic := 'U';
          N_124                : in    std_logic := 'U';
          sFull_RNI9VRD_0      : in    std_logic := 'U';
          N_146                : in    std_logic := 'U';
          N_70                 : in    std_logic := 'U';
          sEmpty_RNI5EFO_0     : in    std_logic := 'U';
          N_33                 : in    std_logic := 'U';
          N_62                 : in    std_logic := 'U';
          N_155                : in    std_logic := 'U';
          sFull_RNI9VRD_1      : in    std_logic := 'U';
          N_147                : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_fifo_ctrlZ6
    port( Waddr_vect_RNI64MA       : out   std_logic_vector(2 to 2);
          data_addr_w_1_iv_i_s_0_0 : in    std_logic_vector(6 to 6) := (others => 'U');
          time_wen                 : in    std_logic_vector(2 to 2) := (others => 'U');
          data_addr_r_0_iv_i_1     : out   std_logic_vector(5 to 5);
          data_addr_r_1_iv_i_s_1   : out   std_logic_vector(6 to 6);
          time_mem_ren_i_0_1       : in    std_logic := 'U';
          data_addr_r_iv_i_a2_0    : out   std_logic_vector(4 to 4);
          data_addr_r_iv_i_1       : out   std_logic_vector(4 downto 0);
          time_ren                 : in    std_logic_vector(2 to 2) := (others => 'U');
          time_ren_1z              : in    std_logic := 'U';
          HRESETn_c                : in    std_logic := 'U';
          HCLK_c                   : in    std_logic := 'U';
          sFull_RNI9VRD_0          : out   std_logic;
          N_147                    : out   std_logic;
          sFull_RNI9VRD_1          : out   std_logic;
          sFull_RNI9VRD            : out   std_logic;
          un13_time_write          : in    std_logic := 'U';
          N_163                    : out   std_logic;
          N_155                    : out   std_logic;
          N_162                    : in    std_logic := 'U';
          sFull_RNIU5GK1           : out   std_logic;
          N_29                     : in    std_logic := 'U';
          N_30_1                   : in    std_logic := 'U';
          N_72                     : in    std_logic := 'U';
          N_56                     : in    std_logic := 'U';
          N_48                     : in    std_logic := 'U';
          N_35                     : in    std_logic := 'U';
          N_64                     : in    std_logic := 'U'
        );
  end component;

    signal N_156, N_89, \time_mem_addr_w_3[0]\, N_132, 
        \time_mem_addr_w_3_i_0[3]\, N_148, \time_mem_addr_w_3[1]\, 
        \data_addr_w_iv_i_2[3]\, \data_addr_w_iv_i_1[3]\, 
        \data_addr_w_iv_i_2[0]\, \data_addr_w_iv_i_1[0]\, 
        \data_addr_w_iv_i_2[1]\, \data_addr_w_iv_i_1[1]\, 
        \Raddr_vect_RNI4A0PH[0]\, \Raddr_vect_RNICA1PH[1]\, 
        \Raddr_vect_RNIKA2PH[2]\, \Raddr_vect_RNIE6Q5I[3]\, 
        \Raddr_vect_RNIIMQ5I[4]\, \Waddr_vect_RNION355[0]\, 
        \Waddr_vect_RNI0O455[1]\, \Waddr_vect_RNI394D5[2]\, 
        \Waddr_vect_RNIJTNE5[3]\, \Waddr_vect_RNILLSP5[4]\, 
        N_1_i_1, sEmpty_RNIE7T87, sEmpty_RNILSD08, sFull_RNIHL443, 
        sFull_RNIU5GK1, N_1_i_1_i, 
        \data_addr_w_1_iv_i_a2_1_1_0[6]\, 
        \data_addr_w_1_iv_i_s_0_0[6]\, \data_mem_ren_i_0[1]\, 
        \time_mem_ren_i_0[3]\, \data_addr_r_1_iv_i_a9_1_1[6]\, 
        N_124, N_64, N_140, N_30_1, N_163, N_164, N_72, N_56, 
        N_48, N_35, N_113, N_162, N_77, \time_mem_ren_i_0[1]\, 
        \data_addr_w_0_iv_i_1[5]\, \Waddr_vect_RNILN58[0]\, 
        \Waddr_vect_RNINV58[2]\, \Waddr_vect_RNI64MA[2]\, 
        \data_addr_w_iv_i_2[2]\, \data_addr_w_iv_i_2[4]\, 
        \time_mem_wen_i_0[0]\, \data_addr_r_0_iv_i_1[5]\, 
        \data_addr_r_0_iv_i_2[5]\, \Raddr_vect_RNI8J9L[2]\, 
        \data_addr_r_iv_i_0[0]\, \data_addr_r_iv_i_0[1]\, 
        \data_addr_r_iv_i_0[2]\, \data_addr_r_iv_i_0[3]\, 
        \data_addr_r_iv_i_0[4]\, sFull_RNI9VRD, sFull_RNIPQBB_0, 
        N_122, sFull_RNI9VRD_0, N_146, N_70, sEmpty_RNI5EFO_0, 
        N_33, N_62, N_155, sFull_RNI9VRD_1, N_147, 
        \data_addr_r_1_iv_i_s_1[6]\, \data_addr_r_iv_i_a2_0[4]\, 
        \data_addr_r_iv_i_1[0]\, \data_addr_r_iv_i_1[1]\, 
        \data_addr_r_iv_i_1[2]\, \data_addr_r_iv_i_1[3]\, 
        \data_addr_r_iv_i_1[4]\, N_29, \data_mem_wen_i_0[2]\, 
        N_128, N_152, N_136, N_68, N_144, N_166, N_160, N_76, 
        N_60, N_52, N_86, N_44, \data_mem_ren_i_0[0]\, 
        \data_mem_wen_i_0[1]\, \data_addr_w_iv_i_4[0]\, 
        \data_addr_w_iv_i_4[1]\, \data_addr_w_iv_i_4[2]\, 
        \data_addr_w_iv_i_4[3]\, \data_addr_w_iv_i_4[4]\, 
        \data_addr_r_iv_i_3[0]\, \data_addr_r_iv_i_3[1]\, 
        \data_addr_r_iv_i_3[2]\, \data_addr_r_iv_i_3[3]\, 
        \data_addr_r_iv_i_3[4]\, N_165, N_120_i, N_158, N_142, 
        N_134, N_126, N_150, \data_addr_r_iv_i_a2_2[4]\, N_67, 
        N_75, N_59, N_51, N_43, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : lpp_waveform_fifo_ctrlZ1
	Use entity work.lpp_waveform_fifo_ctrlZ1(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ7
	Use entity work.lpp_waveform_fifo_ctrlZ7(DEF_ARCH);
    for all : syncram_2pZ1
	Use entity work.syncram_2pZ1(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ2
	Use entity work.lpp_waveform_fifo_ctrlZ2(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ5
	Use entity work.lpp_waveform_fifo_ctrlZ5(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ3
	Use entity work.lpp_waveform_fifo_ctrlZ3(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ0
	Use entity work.lpp_waveform_fifo_ctrlZ0(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ4
	Use entity work.lpp_waveform_fifo_ctrlZ4(DEF_ARCH);
    for all : lpp_waveform_fifo_ctrlZ6
	Use entity work.lpp_waveform_fifo_ctrlZ6(DEF_ARCH);
begin 


    \gen_fifo_ctrl_data.1.lpp_waveform_fifo_ctrl_data\ : 
        lpp_waveform_fifo_ctrlZ1
      port map(ready_i_0(1) => ready_i_0(1), 
        Raddr_vect_RNICA1PH(1) => \Raddr_vect_RNICA1PH[1]\, 
        data_mem_wen_i_0(2) => \data_mem_wen_i_0[2]\, 
        data_mem_wen_i_0(1) => \data_mem_wen_i_0[1]\, 
        Raddr_vect_RNIIMQ5I(4) => \Raddr_vect_RNIIMQ5I[4]\, 
        Raddr_vect_RNIE6Q5I(3) => \Raddr_vect_RNIE6Q5I[3]\, 
        Raddr_vect_RNIKA2PH(2) => \Raddr_vect_RNIKA2PH[2]\, 
        data_addr_r_iv_i_3(4) => \data_addr_r_iv_i_3[4]\, 
        data_addr_r_iv_i_3(3) => \data_addr_r_iv_i_3[3]\, 
        data_addr_r_iv_i_3(2) => \data_addr_r_iv_i_3[2]\, 
        data_addr_r_iv_i_3(1) => \data_addr_r_iv_i_3[1]\, 
        data_addr_r_iv_i_3(0) => \data_addr_r_iv_i_3[0]\, 
        Raddr_vect_RNI4A0PH(0) => \Raddr_vect_RNI4A0PH[0]\, 
        data_addr_r_iv_i_a2_2(4) => \data_addr_r_iv_i_a2_2[4]\, 
        data_wen(1) => data_wen(1), data_mem_ren_i_0(1) => 
        \data_mem_ren_i_0[1]\, data_mem_ren_i_0(0) => 
        \data_mem_ren_i_0[0]\, data_ren(1) => data_ren(1), 
        data_ren_1z => data_ren_1z, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, N_166 => N_166, N_126 => N_126, N_150
         => N_150, N_134 => N_134, N_142 => N_142, N_165 => N_165, 
        N_158 => N_158, un20_time_write => un20_time_write, N_68
         => N_68, N_164 => N_164, N_120_i => N_120_i, N_44 => 
        N_44, N_52 => N_52, N_60 => N_60, N_76 => N_76, N_86 => 
        N_86, N_75 => N_75, N_59 => N_59, N_51 => N_51, N_43 => 
        N_43, N_67 => N_67);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \gen_fifo_ctrl_time.3.lpp_waveform_fifo_ctrl_time\ : 
        lpp_waveform_fifo_ctrlZ7
      port map(time_mem_addr_w_3_i_0_1 => 
        \time_mem_addr_w_3_i_0[3]\, 
        data_addr_w_1_iv_i_a2_1_1_0(6) => 
        \data_addr_w_1_iv_i_a2_1_1_0[6]\, 
        data_addr_w_1_iv_i_s_0_0(6) => 
        \data_addr_w_1_iv_i_s_0_0[6]\, time_wen(3) => time_wen(3), 
        time_ren(3) => time_ren(3), data_mem_ren_i_0(1) => 
        \data_mem_ren_i_0[1]\, time_mem_ren_i_0(3) => 
        \time_mem_ren_i_0[3]\, data_addr_r_1_iv_i_a9_1_1(6) => 
        \data_addr_r_1_iv_i_a9_1_1[6]\, time_mem_addr_w_3(1) => 
        \time_mem_addr_w_3[1]\, time_mem_addr_w_3(0) => 
        \time_mem_addr_w_3[0]\, HRESETn_c => HRESETn_c, HCLK_c
         => HCLK_c, N_124 => N_124, N_64 => N_64, N_140 => N_140, 
        N_30_1 => N_30_1, N_89 => N_89, N_163 => N_163, N_164 => 
        N_164, N_72 => N_72, N_56 => N_56, N_48 => N_48, N_35 => 
        N_35, N_113 => N_113, N_162 => N_162, N_77 => N_77);
    
    SRAM : syncram_2pZ1
      port map(hwdata_c(31) => hwdata_c(31), hwdata_c(30) => 
        hwdata_c(30), hwdata_c(29) => hwdata_c(29), hwdata_c(28)
         => hwdata_c(28), hwdata_c(27) => hwdata_c(27), 
        hwdata_c(26) => hwdata_c(26), hwdata_c(25) => 
        hwdata_c(25), hwdata_c(24) => hwdata_c(24), hwdata_c(23)
         => hwdata_c(23), hwdata_c(22) => hwdata_c(22), 
        hwdata_c(21) => hwdata_c(21), hwdata_c(20) => 
        hwdata_c(20), hwdata_c(19) => hwdata_c(19), hwdata_c(18)
         => hwdata_c(18), hwdata_c(17) => hwdata_c(17), 
        hwdata_c(16) => hwdata_c(16), hwdata_c(15) => 
        hwdata_c(15), hwdata_c(14) => hwdata_c(14), hwdata_c(13)
         => hwdata_c(13), hwdata_c(12) => hwdata_c(12), 
        hwdata_c(11) => hwdata_c(11), hwdata_c(10) => 
        hwdata_c(10), hwdata_c(9) => hwdata_c(9), hwdata_c(8) => 
        hwdata_c(8), hwdata_c(7) => hwdata_c(7), hwdata_c(6) => 
        hwdata_c(6), hwdata_c(5) => hwdata_c(5), hwdata_c(4) => 
        hwdata_c(4), hwdata_c(3) => hwdata_c(3), hwdata_c(2) => 
        hwdata_c(2), hwdata_c(1) => hwdata_c(1), hwdata_c(0) => 
        hwdata_c(0), Raddr_vect_RNI4A0PH(0) => 
        \Raddr_vect_RNI4A0PH[0]\, Raddr_vect_RNICA1PH(1) => 
        \Raddr_vect_RNICA1PH[1]\, Raddr_vect_RNIKA2PH(2) => 
        \Raddr_vect_RNIKA2PH[2]\, Raddr_vect_RNIE6Q5I(3) => 
        \Raddr_vect_RNIE6Q5I[3]\, Raddr_vect_RNIIMQ5I(4) => 
        \Raddr_vect_RNIIMQ5I[4]\, Waddr_vect_RNION355(0) => 
        \Waddr_vect_RNION355[0]\, Waddr_vect_RNI0O455(1) => 
        \Waddr_vect_RNI0O455[1]\, Waddr_vect_RNI394D5(2) => 
        \Waddr_vect_RNI394D5[2]\, Waddr_vect_RNIJTNE5(3) => 
        \Waddr_vect_RNIJTNE5[3]\, Waddr_vect_RNILLSP5(4) => 
        \Waddr_vect_RNILLSP5[4]\, wdata(31) => wdata(31), 
        wdata(30) => wdata(30), wdata(29) => wdata(29), wdata(28)
         => wdata(28), wdata(27) => wdata(27), wdata(26) => 
        wdata(26), wdata(25) => wdata(25), wdata(24) => wdata(24), 
        wdata(23) => wdata(23), wdata(22) => wdata(22), wdata(21)
         => wdata(21), wdata(20) => wdata(20), wdata(19) => 
        wdata(19), wdata(18) => wdata(18), wdata(17) => wdata(17), 
        wdata(16) => wdata(16), wdata(15) => wdata(15), wdata(14)
         => wdata(14), wdata(13) => wdata(13), wdata(12) => 
        wdata(12), wdata(11) => wdata(11), wdata(10) => wdata(10), 
        wdata(9) => wdata(9), wdata(8) => wdata(8), wdata(7) => 
        wdata(7), wdata(6) => wdata(6), wdata(5) => wdata(5), 
        wdata(4) => wdata(4), wdata(3) => wdata(3), wdata(2) => 
        wdata(2), wdata(1) => wdata(1), wdata(0) => wdata(0), 
        HCLK_c => HCLK_c, N_1_i_1 => N_1_i_1, sEmpty_RNIE7T87 => 
        sEmpty_RNIE7T87, sEmpty_RNILSD08 => sEmpty_RNILSD08, 
        sFull_RNIHL443 => sFull_RNIHL443, sFull_RNIU5GK1 => 
        sFull_RNIU5GK1, syncram_2pZ1_GND => lpp_waveform_fifo_GND, 
        syncram_2pZ1_VCC => lpp_waveform_fifo_VCC, N_1_i_1_i => 
        N_1_i_1_i);
    
    \data_addr_w_iv_i_a2_2[0]\ : OR2A
      port map(A => N_89, B => \time_mem_addr_w_3[0]\, Y => N_156);
    
    \data_addr_w_iv_i_a2_2_RNIRMOT[0]\ : AND2
      port map(A => \data_addr_w_iv_i_1[0]\, B => N_156, Y => 
        \data_addr_w_iv_i_2[0]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \gen_fifo_ctrl_data.2.lpp_waveform_fifo_ctrl_data\ : 
        lpp_waveform_fifo_ctrlZ2
      port map(ready_i_0(2) => ready_i_0(2), data_mem_wen_i_0(2)
         => \data_mem_wen_i_0[2]\, data_ren(2) => data_ren(2), 
        Waddr_vect_RNI0O455(1) => \Waddr_vect_RNI0O455[1]\, 
        Waddr_vect_RNILLSP5(4) => \Waddr_vect_RNILLSP5[4]\, 
        Waddr_vect_RNIJTNE5(3) => \Waddr_vect_RNIJTNE5[3]\, 
        Waddr_vect_RNI394D5(2) => \Waddr_vect_RNI394D5[2]\, 
        data_mem_ren_i_0_0 => \data_mem_ren_i_0[0]\, 
        data_addr_r_0_iv_i_2(5) => \data_addr_r_0_iv_i_2[5]\, 
        data_addr_w_iv_i_4(4) => \data_addr_w_iv_i_4[4]\, 
        data_addr_w_iv_i_4(3) => \data_addr_w_iv_i_4[3]\, 
        data_addr_w_iv_i_4(2) => \data_addr_w_iv_i_4[2]\, 
        data_addr_w_iv_i_4(1) => \data_addr_w_iv_i_4[1]\, 
        data_addr_w_iv_i_4(0) => \data_addr_w_iv_i_4[0]\, 
        Waddr_vect_RNION355(0) => \Waddr_vect_RNION355[0]\, 
        data_wen(2) => data_wen(2), data_addr_r_iv_i_a2_0(4) => 
        \data_addr_r_iv_i_a2_0[4]\, data_addr_r_iv_i_a2_2(4) => 
        \data_addr_r_iv_i_a2_2[4]\, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, N_67 => N_67, N_166 => N_166, N_75 => 
        N_75, N_59 => N_59, N_51 => N_51, N_43 => N_43, N_152 => 
        N_152, N_128 => N_128, N_136 => N_136, N_144 => N_144, 
        sEmpty_RNIE7T87 => sEmpty_RNIE7T87, N_160 => N_160, N_77
         => N_77);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \gen_fifo_ctrl_time.1.lpp_waveform_fifo_ctrl_time\ : 
        lpp_waveform_fifo_ctrlZ5
      port map(time_mem_wen_i_0_0 => \time_mem_wen_i_0[0]\, 
        Waddr_vect_RNINV58(2) => \Waddr_vect_RNINV58[2]\, 
        Waddr_vect_RNILN58(0) => \Waddr_vect_RNILN58[0]\, 
        Raddr_vect_RNI8J9L(2) => \Raddr_vect_RNI8J9L[2]\, 
        time_mem_ren_i_0(1) => \time_mem_ren_i_0[1]\, time_wen(1)
         => time_wen(1), time_ren(1) => time_ren(1), HRESETn_c
         => HRESETn_c, HCLK_c => HCLK_c, N_146 => N_146, N_162
         => N_162, N_113 => N_113, N_122 => N_122, 
        sFull_RNIPQBB_0 => sFull_RNIPQBB_0, N_62 => N_62, N_70
         => N_70, sEmpty_RNI5EFO_0 => sEmpty_RNI5EFO_0, N_33 => 
        N_33, N_29 => N_29);
    
    \gen_fifo_ctrl_data.3.lpp_waveform_fifo_ctrl_data\ : 
        lpp_waveform_fifo_ctrlZ3
      port map(ready_i_0(3) => ready_i_0(3), data_mem_wen_i_0_0
         => \data_mem_wen_i_0[2]\, data_ren(3) => data_ren(3), 
        data_wen(3) => data_wen(3), HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, N_128 => N_128, N_152 => N_152, N_136
         => N_136, N_68 => N_68, N_144 => N_144, N_166 => N_166, 
        N_160 => N_160, N_76 => N_76, N_60 => N_60, N_52 => N_52, 
        N_86 => N_86, N_44 => N_44, N_1_i_1 => N_1_i_1, N_1_i_1_i
         => N_1_i_1_i);
    
    \gen_fifo_ctrl_data.0.lpp_waveform_fifo_ctrl_data\ : 
        lpp_waveform_fifo_ctrlZ0
      port map(ready_i_0(0) => ready_i_0(0), data_ren(0) => 
        data_ren(0), data_addr_w_0_iv_i_1(5) => 
        \data_addr_w_0_iv_i_1[5]\, data_addr_r_1_iv_i_s_1(6) => 
        \data_addr_r_1_iv_i_s_1[6]\, data_addr_r_1_iv_i_a9_1_1(6)
         => \data_addr_r_1_iv_i_a9_1_1[6]\, data_mem_ren_i_0(0)
         => \data_mem_ren_i_0[0]\, data_mem_wen_i_0_1 => 
        \data_mem_wen_i_0[1]\, data_addr_w_1_iv_i_a2_1_1_0(6) => 
        \data_addr_w_1_iv_i_a2_1_1_0[6]\, data_addr_w_iv_i_2(4)
         => \data_addr_w_iv_i_2[4]\, data_addr_w_iv_i_2(3) => 
        \data_addr_w_iv_i_2[3]\, data_addr_w_iv_i_2(2) => 
        \data_addr_w_iv_i_2[2]\, data_addr_w_iv_i_2(1) => 
        \data_addr_w_iv_i_2[1]\, data_addr_w_iv_i_2(0) => 
        \data_addr_w_iv_i_2[0]\, data_addr_w_iv_i_4(4) => 
        \data_addr_w_iv_i_4[4]\, data_addr_w_iv_i_4(3) => 
        \data_addr_w_iv_i_4[3]\, data_addr_w_iv_i_4(2) => 
        \data_addr_w_iv_i_4[2]\, data_addr_w_iv_i_4(1) => 
        \data_addr_w_iv_i_4[1]\, data_addr_w_iv_i_4(0) => 
        \data_addr_w_iv_i_4[0]\, data_wen(0) => data_wen(0), 
        data_addr_r_iv_i_0(4) => \data_addr_r_iv_i_0[4]\, 
        data_addr_r_iv_i_0(3) => \data_addr_r_iv_i_0[3]\, 
        data_addr_r_iv_i_0(2) => \data_addr_r_iv_i_0[2]\, 
        data_addr_r_iv_i_0(1) => \data_addr_r_iv_i_0[1]\, 
        data_addr_r_iv_i_0(0) => \data_addr_r_iv_i_0[0]\, 
        data_addr_r_iv_i_1(4) => \data_addr_r_iv_i_1[4]\, 
        data_addr_r_iv_i_1(3) => \data_addr_r_iv_i_1[3]\, 
        data_addr_r_iv_i_1(2) => \data_addr_r_iv_i_1[2]\, 
        data_addr_r_iv_i_1(1) => \data_addr_r_iv_i_1[1]\, 
        data_addr_r_iv_i_1(0) => \data_addr_r_iv_i_1[0]\, 
        data_addr_r_iv_i_3(4) => \data_addr_r_iv_i_3[4]\, 
        data_addr_r_iv_i_3(3) => \data_addr_r_iv_i_3[3]\, 
        data_addr_r_iv_i_3(2) => \data_addr_r_iv_i_3[2]\, 
        data_addr_r_iv_i_3(1) => \data_addr_r_iv_i_3[1]\, 
        data_addr_r_iv_i_3(0) => \data_addr_r_iv_i_3[0]\, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, N_165 => N_165, 
        N_120_i => N_120_i, sFull_RNIHL443 => sFull_RNIHL443, 
        sEmpty_RNILSD08 => sEmpty_RNILSD08, N_124 => N_124, N_164
         => N_164, N_158 => N_158, N_142 => N_142, N_134 => N_134, 
        N_126 => N_126, N_150 => N_150);
    
    \data_addr_w_iv_i_a2_2_RNIACB71[3]\ : AND2
      port map(A => N_132, B => \data_addr_w_iv_i_1[3]\, Y => 
        \data_addr_w_iv_i_2[3]\);
    
    \data_addr_w_iv_i_a2_2[3]\ : NAND2
      port map(A => N_89, B => \time_mem_addr_w_3_i_0[3]\, Y => 
        N_132);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \gen_fifo_ctrl_time.0.lpp_waveform_fifo_ctrl_time\ : 
        lpp_waveform_fifo_ctrlZ4
      port map(time_mem_ren_i_0_1 => \time_mem_ren_i_0[1]\, 
        time_wen(0) => time_wen(0), time_ren(0) => time_ren(0), 
        data_addr_w_0_iv_i_1(5) => \data_addr_w_0_iv_i_1[5]\, 
        Waddr_vect_RNILN58(0) => \Waddr_vect_RNILN58[0]\, 
        Waddr_vect_RNINV58(2) => \Waddr_vect_RNINV58[2]\, 
        Waddr_vect_RNI64MA(2) => \Waddr_vect_RNI64MA[2]\, 
        data_addr_w_iv_i_2_0 => \data_addr_w_iv_i_2[2]\, 
        data_addr_w_iv_i_2_2 => \data_addr_w_iv_i_2[4]\, 
        time_mem_wen_i_0(0) => \time_mem_wen_i_0[0]\, 
        data_addr_r_0_iv_i_1(5) => \data_addr_r_0_iv_i_1[5]\, 
        data_addr_r_0_iv_i_2(5) => \data_addr_r_0_iv_i_2[5]\, 
        Raddr_vect_RNI8J9L(2) => \Raddr_vect_RNI8J9L[2]\, 
        data_addr_r_iv_i_0(4) => \data_addr_r_iv_i_0[4]\, 
        data_addr_r_iv_i_0(3) => \data_addr_r_iv_i_0[3]\, 
        data_addr_r_iv_i_0(2) => \data_addr_r_iv_i_0[2]\, 
        data_addr_r_iv_i_0(1) => \data_addr_r_iv_i_0[1]\, 
        data_addr_r_iv_i_0(0) => \data_addr_r_iv_i_0[0]\, 
        data_addr_w_iv_i_1_0 => \data_addr_w_iv_i_1[0]\, 
        data_addr_w_iv_i_1_3 => \data_addr_w_iv_i_1[3]\, 
        data_addr_w_iv_i_1_1 => \data_addr_w_iv_i_1[1]\, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, N_77 => N_77, 
        sFull_RNI9VRD => sFull_RNI9VRD, N_140 => N_140, 
        sFull_RNIPQBB_0 => sFull_RNIPQBB_0, N_122 => N_122, N_124
         => N_124, sFull_RNI9VRD_0 => sFull_RNI9VRD_0, N_146 => 
        N_146, N_70 => N_70, sEmpty_RNI5EFO_0 => sEmpty_RNI5EFO_0, 
        N_33 => N_33, N_62 => N_62, N_155 => N_155, 
        sFull_RNI9VRD_1 => sFull_RNI9VRD_1, N_147 => N_147);
    
    \data_addr_w_iv_i_a2_2[1]\ : OR2A
      port map(A => N_89, B => \time_mem_addr_w_3[1]\, Y => N_148);
    
    \gen_fifo_ctrl_time.2.lpp_waveform_fifo_ctrl_time\ : 
        lpp_waveform_fifo_ctrlZ6
      port map(Waddr_vect_RNI64MA(2) => \Waddr_vect_RNI64MA[2]\, 
        data_addr_w_1_iv_i_s_0_0(6) => 
        \data_addr_w_1_iv_i_s_0_0[6]\, time_wen(2) => time_wen(2), 
        data_addr_r_0_iv_i_1(5) => \data_addr_r_0_iv_i_1[5]\, 
        data_addr_r_1_iv_i_s_1(6) => \data_addr_r_1_iv_i_s_1[6]\, 
        time_mem_ren_i_0_1 => \time_mem_ren_i_0[3]\, 
        data_addr_r_iv_i_a2_0(4) => \data_addr_r_iv_i_a2_0[4]\, 
        data_addr_r_iv_i_1(4) => \data_addr_r_iv_i_1[4]\, 
        data_addr_r_iv_i_1(3) => \data_addr_r_iv_i_1[3]\, 
        data_addr_r_iv_i_1(2) => \data_addr_r_iv_i_1[2]\, 
        data_addr_r_iv_i_1(1) => \data_addr_r_iv_i_1[1]\, 
        data_addr_r_iv_i_1(0) => \data_addr_r_iv_i_1[0]\, 
        time_ren(2) => time_ren(2), time_ren_1z => time_ren_1z, 
        HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, sFull_RNI9VRD_0
         => sFull_RNI9VRD_0, N_147 => N_147, sFull_RNI9VRD_1 => 
        sFull_RNI9VRD_1, sFull_RNI9VRD => sFull_RNI9VRD, 
        un13_time_write => un13_time_write, N_163 => N_163, N_155
         => N_155, N_162 => N_162, sFull_RNIU5GK1 => 
        sFull_RNIU5GK1, N_29 => N_29, N_30_1 => N_30_1, N_72 => 
        N_72, N_56 => N_56, N_48 => N_48, N_35 => N_35, N_64 => 
        N_64);
    
    \data_addr_w_iv_i_a2_2_RNIV6PT[1]\ : AND2
      port map(A => \data_addr_w_iv_i_1[1]\, B => N_148, Y => 
        \data_addr_w_iv_i_2[1]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_snapshot_160_11 is

    port( sample_f0_wdata_95 : in    std_logic;
          sample_f0_wdata_94 : in    std_logic;
          sample_f0_wdata_93 : in    std_logic;
          sample_f0_wdata_92 : in    std_logic;
          sample_f0_wdata_91 : in    std_logic;
          sample_f0_wdata_90 : in    std_logic;
          sample_f0_wdata_89 : in    std_logic;
          sample_f0_wdata_88 : in    std_logic;
          sample_f0_wdata_87 : in    std_logic;
          sample_f0_wdata_86 : in    std_logic;
          sample_f0_wdata_85 : in    std_logic;
          sample_f0_wdata_84 : in    std_logic;
          sample_f0_wdata_83 : in    std_logic;
          sample_f0_wdata_82 : in    std_logic;
          sample_f0_wdata_81 : in    std_logic;
          sample_f0_wdata_80 : in    std_logic;
          sample_f0_wdata_79 : in    std_logic;
          sample_f0_wdata_78 : in    std_logic;
          sample_f0_wdata_77 : in    std_logic;
          sample_f0_wdata_76 : in    std_logic;
          sample_f0_wdata_75 : in    std_logic;
          sample_f0_wdata_74 : in    std_logic;
          sample_f0_wdata_73 : in    std_logic;
          sample_f0_wdata_72 : in    std_logic;
          sample_f0_wdata_71 : in    std_logic;
          sample_f0_wdata_70 : in    std_logic;
          sample_f0_wdata_69 : in    std_logic;
          sample_f0_wdata_68 : in    std_logic;
          sample_f0_wdata_67 : in    std_logic;
          sample_f0_wdata_66 : in    std_logic;
          sample_f0_wdata_65 : in    std_logic;
          sample_f0_wdata_64 : in    std_logic;
          sample_f0_wdata_63 : in    std_logic;
          sample_f0_wdata_62 : in    std_logic;
          sample_f0_wdata_61 : in    std_logic;
          sample_f0_wdata_60 : in    std_logic;
          sample_f0_wdata_59 : in    std_logic;
          sample_f0_wdata_58 : in    std_logic;
          sample_f0_wdata_57 : in    std_logic;
          sample_f0_wdata_56 : in    std_logic;
          sample_f0_wdata_55 : in    std_logic;
          sample_f0_wdata_54 : in    std_logic;
          sample_f0_wdata_53 : in    std_logic;
          sample_f0_wdata_52 : in    std_logic;
          sample_f0_wdata_51 : in    std_logic;
          sample_f0_wdata_50 : in    std_logic;
          sample_f0_wdata_49 : in    std_logic;
          sample_f0_wdata_48 : in    std_logic;
          sample_f0_wdata_15 : in    std_logic;
          sample_f0_wdata_14 : in    std_logic;
          sample_f0_wdata_13 : in    std_logic;
          sample_f0_wdata_12 : in    std_logic;
          sample_f0_wdata_11 : in    std_logic;
          sample_f0_wdata_10 : in    std_logic;
          sample_f0_wdata_9  : in    std_logic;
          sample_f0_wdata_8  : in    std_logic;
          sample_f0_wdata_7  : in    std_logic;
          sample_f0_wdata_6  : in    std_logic;
          sample_f0_wdata_5  : in    std_logic;
          sample_f0_wdata_4  : in    std_logic;
          sample_f0_wdata_3  : in    std_logic;
          sample_f0_wdata_2  : in    std_logic;
          sample_f0_wdata_1  : in    std_logic;
          sample_f0_wdata_0  : in    std_logic;
          data_f0_out        : out   std_logic_vector(159 downto 64);
          nb_snapshot_param  : in    std_logic_vector(10 downto 0);
          sample_f0_37       : in    std_logic;
          sample_f0_5        : in    std_logic;
          sample_f0_38       : in    std_logic;
          sample_f0_6        : in    std_logic;
          sample_f0_39       : in    std_logic;
          sample_f0_7        : in    std_logic;
          sample_f0_40       : in    std_logic;
          sample_f0_8        : in    std_logic;
          sample_f0_41       : in    std_logic;
          sample_f0_9        : in    std_logic;
          sample_f0_42       : in    std_logic;
          sample_f0_10       : in    std_logic;
          sample_f0_43       : in    std_logic;
          sample_f0_11       : in    std_logic;
          sample_f0_61       : in    std_logic;
          sample_f0_62       : in    std_logic;
          sample_f0_63       : in    std_logic;
          sample_f0_32       : in    std_logic;
          sample_f0_0        : in    std_logic;
          sample_f0_33       : in    std_logic;
          sample_f0_1        : in    std_logic;
          sample_f0_34       : in    std_logic;
          sample_f0_2        : in    std_logic;
          sample_f0_35       : in    std_logic;
          sample_f0_3        : in    std_logic;
          sample_f0_36       : in    std_logic;
          sample_f0_4        : in    std_logic;
          sample_f0_48       : in    std_logic;
          sample_f0_49       : in    std_logic;
          sample_f0_50       : in    std_logic;
          sample_f0_51       : in    std_logic;
          sample_f0_52       : in    std_logic;
          sample_f0_53       : in    std_logic;
          sample_f0_54       : in    std_logic;
          sample_f0_55       : in    std_logic;
          sample_f0_56       : in    std_logic;
          sample_f0_57       : in    std_logic;
          sample_f0_58       : in    std_logic;
          sample_f0_59       : in    std_logic;
          sample_f0_60       : in    std_logic;
          sample_f0_44       : in    std_logic;
          sample_f0_12       : in    std_logic;
          sample_f0_45       : in    std_logic;
          sample_f0_13       : in    std_logic;
          sample_f0_46       : in    std_logic;
          sample_f0_14       : in    std_logic;
          sample_f0_47       : in    std_logic;
          sample_f0_15       : in    std_logic;
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic;
          data_f0_out_valid  : out   std_logic;
          enable_f0          : in    std_logic;
          data_shaping_R0    : in    std_logic;
          data_shaping_R0_0  : in    std_logic;
          start_snapshot_f0  : in    std_logic;
          sample_f0_val_0    : in    std_logic;
          burst_f0           : in    std_logic
        );

end lpp_waveform_snapshot_160_11;

architecture DEF_ARCH of lpp_waveform_snapshot_160_11 is 

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \un1_data_out_valid_0_sqmuxa_1_1[31]\, 
        data_out_valid_0_sqmuxa_1, 
        \counter_points_snapshot_0_sqmuxa_1_0\, 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, 
        \data_out_valid_0_sqmuxa\, ADD_32x32_fast_I311_Y_0_0, 
        \counter_points_snapshot[31]_net_1\, 
        ADD_32x32_fast_I308_Y_0_0, 
        \un1_counter_points_snapshot[3]\, 
        ADD_32x32_fast_I296_Y_0_0, 
        \un1_counter_points_snapshot[15]\, 
        ADD_32x32_fast_I310_Y_0_0, 
        \counter_points_snapshot[30]_net_1\, 
        ADD_32x32_fast_I250_Y_2, ADD_32x32_fast_I250_Y_1, N483, 
        N487, N467, N470, N479, ADD_32x32_fast_I304_Y_0_0, 
        \un1_counter_points_snapshot[7]\, 
        ADD_32x32_fast_I253_Y_0_0, I94_un1_Y, N485, 
        ADD_32x32_fast_I295_Y_0_0, 
        \un1_counter_points_snapshot[16]\, 
        ADD_32x32_fast_I303_Y_0_0, 
        \un1_counter_points_snapshot[8]\, 
        ADD_32x32_fast_I288_Y_0_0, 
        \un1_counter_points_snapshot[23]\, 
        ADD_32x32_fast_I251_Y_2, ADD_32x32_fast_I251_Y_1, N489, 
        N464, ADD_32x32_fast_I302_Y_0_0, 
        \un1_counter_points_snapshot[9]\, 
        ADD_32x32_fast_I307_Y_0_0, 
        \un1_counter_points_snapshot[4]\, 
        ADD_32x32_fast_I294_Y_0_0, 
        \un1_counter_points_snapshot[17]\, 
        ADD_32x32_fast_I292_Y_0_0, 
        \un1_counter_points_snapshot[19]\, 
        ADD_32x32_fast_I309_Y_0_0, 
        \counter_points_snapshot[29]_net_1\, 
        ADD_32x32_fast_I300_Y_0_0, 
        \un1_counter_points_snapshot[11]\, 
        ADD_32x32_fast_I306_Y_0_0, 
        \un1_counter_points_snapshot[5]\, 
        ADD_32x32_fast_I305_Y_0_0, 
        \un1_counter_points_snapshot[6]\, 
        ADD_32x32_fast_I287_Y_0_0, 
        \un1_counter_points_snapshot[24]\, 
        ADD_32x32_fast_I291_Y_0_0, 
        \un1_counter_points_snapshot[20]\, 
        ADD_32x32_fast_I299_Y_0_0, 
        \un1_counter_points_snapshot[12]\, 
        ADD_32x32_fast_I301_Y_0_0, 
        \un1_counter_points_snapshot[10]\, 
        ADD_32x32_fast_I254_Y_0, N554, ADD_32x32_fast_I259_Y_0, 
        N636, N620, ADD_32x32_fast_I297_Y_0_0, 
        \counter_points_snapshot[17]_net_1\, 
        ADD_32x32_fast_I298_Y_0_0, 
        \un1_counter_points_snapshot[13]\, 
        ADD_32x32_fast_I252_Y_1, ADD_32x32_fast_I252_Y_0, N491, 
        ADD_32x32_fast_I289_Y_0_0, 
        \un1_counter_points_snapshot[22]\, 
        ADD_32x32_fast_I255_Y_0, N556, ADD_32x32_fast_I293_Y_0_0, 
        \un1_counter_points_snapshot[18]\, 
        ADD_32x32_fast_I256_Y_0, N558, ADD_32x32_fast_I284_Y_0_0, 
        \un1_counter_points_snapshot[27]\, 
        ADD_32x32_fast_I263_Y_0, N644, N628, 
        ADD_32x32_fast_I283_Y_0_0, 
        \un1_counter_points_snapshot[28]\, 
        ADD_32x32_fast_I142_Y_0, 
        \un1_counter_points_snapshot[26]\, 
        ADD_32x32_fast_I118_Y_0, ADD_32x32_fast_I110_Y_0, 
        ADD_32x32_fast_I134_Y_0, 
        \un1_counter_points_snapshot[25]\, 
        ADD_32x32_fast_I126_Y_1, 
        \un1_counter_points_snapshot[21]\, 
        data_out_valid_0_sqmuxa_1_1, un4_data_in_validlt30_27, 
        un4_data_in_validlt30_18, un4_data_in_validlt30_17, 
        un4_data_in_validlt30_23, un4_data_in_validlt30_26, 
        un4_data_in_validlt30_12, un4_data_in_validlt30_11, 
        un4_data_in_validlt30_22, un4_data_in_validlt30_25, 
        un4_data_in_validlt30_8, un4_data_in_validlt30_7, 
        un4_data_in_validlt30_20, un4_data_in_validlt30_2, 
        un4_data_in_validlt30_1, un4_data_in_validlt30_15, 
        un4_data_in_validlt30_14, 
        \counter_points_snapshot[27]_net_1\, 
        \counter_points_snapshot[26]_net_1\, 
        un4_data_in_validlt30_10, 
        \counter_points_snapshot[19]_net_1\, 
        \counter_points_snapshot[18]_net_1\, 
        un4_data_in_validlt30_6, 
        \counter_points_snapshot[11]_net_1\, 
        \counter_points_snapshot[10]_net_1\, 
        un4_data_in_validlt30_4, 
        \counter_points_snapshot[7]_net_1\, 
        \counter_points_snapshot[6]_net_1\, 
        \counter_points_snapshot[1]_net_1\, 
        \counter_points_snapshot[0]_net_1\, 
        \counter_points_snapshot[28]_net_1\, 
        \counter_points_snapshot[24]_net_1\, 
        \counter_points_snapshot[25]_net_1\, 
        \counter_points_snapshot[22]_net_1\, 
        \counter_points_snapshot[23]_net_1\, 
        \counter_points_snapshot[20]_net_1\, 
        \counter_points_snapshot[21]_net_1\, 
        \counter_points_snapshot[16]_net_1\, 
        \counter_points_snapshot[14]_net_1\, 
        \counter_points_snapshot[15]_net_1\, 
        \counter_points_snapshot[12]_net_1\, 
        \counter_points_snapshot[13]_net_1\, 
        \counter_points_snapshot[8]_net_1\, 
        \counter_points_snapshot[9]_net_1\, 
        \counter_points_snapshot[4]_net_1\, 
        \counter_points_snapshot[5]_net_1\, 
        \counter_points_snapshot[2]_net_1\, 
        \counter_points_snapshot[3]_net_1\, 
        \un1_data_out_valid_0_sqmuxa_2[4]\, N533, N529, N754, 
        N634, N618, N650, un4_data_in_validlto30_i, N740, N774, 
        N764, N738, N771, N744, N752, 
        \un1_data_out_valid_0_sqmuxa_2[6]\, N652_i, 
        \un1_data_out_valid_0_sqmuxa_2[1]\, 
        \un1_counter_points_snapshot[30]\, N380, 
        \un1_data_out_valid_0_sqmuxa_2[2]\, 
        \un1_counter_points_snapshot[29]\, 
        \un1_data_out_valid_0_sqmuxa_2[5]\, N654, 
        \un1_data_out_valid_0_sqmuxa_2[8]\, N401, 
        \un1_data_out_valid_0_sqmuxa_2[10]\, N786, N750, N630, 
        N789, \un1_data_out_valid_0_sqmuxa_2[9]\, N756, N748, 
        N497, N766, N646, N746, N626, N783, N572, N419, I66_un1_Y, 
        N580, N407, N588, \un1_data_out_valid_0_sqmuxa_2[3]\, 
        N594, \un1_data_out_valid_0_sqmuxa_2[7]\, N762, N642, 
        N564, I60_un1_Y, N431, N758, N622, N638, N742, N777, 
        \sample_f0_wdata[32]\, \sample_f0_wdata[33]\, 
        \sample_f0_wdata[34]\, \sample_f0_wdata[35]\, 
        \sample_f0_wdata[19]\, \sample_f0_wdata[20]\, 
        \sample_f0_wdata[21]\, \sample_f0_wdata[22]\, 
        \sample_f0_wdata[23]\, \sample_f0_wdata[24]\, 
        \sample_f0_wdata[25]\, \sample_f0_wdata[26]\, 
        \sample_f0_wdata[27]\, \sample_f0_wdata[28]\, 
        \sample_f0_wdata[29]\, \sample_f0_wdata[30]\, 
        \sample_f0_wdata[31]\, \sample_f0_wdata[43]\, 
        \sample_f0_wdata[44]\, \sample_f0_wdata[45]\, 
        \sample_f0_wdata[46]\, \sample_f0_wdata[47]\, 
        \sample_f0_wdata[16]\, \sample_f0_wdata[17]\, 
        \sample_f0_wdata[18]\, \sample_f0_wdata[36]\, 
        \sample_f0_wdata[37]\, \sample_f0_wdata[38]\, 
        \sample_f0_wdata[39]\, \sample_f0_wdata[40]\, 
        \sample_f0_wdata[41]\, \sample_f0_wdata[42]\, 
        \counter_points_snapshot_10[4]\, N_90, 
        \counter_points_snapshot_2_sqmuxa\, 
        \counter_points_snapshot_10[23]\, 
        un1_counter_points_snapshot_0_sqmuxa_1_i, N461, 
        \counter_points_snapshot_3_sqmuxa\, 
        \un1_data_out_valid_0_sqmuxa_1[31]\, 
        counter_points_snapshot_0_sqmuxa_i, data_out_valid_19, 
        un1_enable_2, \counter_points_snapshot_10[30]\, 
        \counter_points_snapshot_0_sqmuxa_1\, 
        \counter_points_snapshot_10[31]\, 
        \counter_points_snapshot_10[22]\, 
        \counter_points_snapshot_10[24]\, 
        \counter_points_snapshot_10[28]\, N760, 
        \counter_points_snapshot_10[18]\, N590, N582, N_92, 
        \counter_points_snapshot_2_sqmuxa_2\, 
        \counter_points_snapshot_10[6]\, N507, N511, N578, N586, 
        I74_un1_Y, \un1_counter_points_snapshot[31]\, 
        \counter_points_snapshot_10[10]\, N_96, 
        \counter_points_snapshot_10[8]\, N_94, 
        \counter_points_snapshot_10[5]\, N_91, 
        \counter_points_snapshot_10[2]\, N_88, 
        \counter_points_snapshot_10[1]\, N_87, N562, 
        \counter_points_snapshot_10[25]\, N_95, 
        \counter_points_snapshot_10[9]\, 
        \counter_points_snapshot_10[27]\, 
        \counter_points_snapshot_10[26]\, 
        \counter_points_snapshot_10[17]\, 
        \counter_points_snapshot_10[14]\, 
        \counter_points_snapshot_10[15]\, 
        \counter_points_snapshot_10[11]\, N515, 
        \counter_points_snapshot_10[16]\, N768, N523, N531, N527, 
        \un1_data_out_valid_0_sqmuxa_2[0]\, N_86, 
        \counter_points_snapshot_10[0]\, 
        \counter_points_snapshot_10[19]\, 
        \counter_points_snapshot_10[7]\, N_93, 
        \counter_points_snapshot_10[3]\, N_89, 
        \counter_points_snapshot_10[20]\, N434, N780, 
        \counter_points_snapshot_10[12]\, 
        \counter_points_snapshot_10[29]\, 
        \counter_points_snapshot_10[21]\, 
        \counter_points_snapshot_10[13]\, N574, N566, N503, N495, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \counter_points_snapshot_RNIV49P[18]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[18]_net_1\, Y => 
        \un1_counter_points_snapshot[13]\);
    
    \counter_points_snapshot_RNIRF66[2]\ : NOR2
      port map(A => \counter_points_snapshot[2]_net_1\, B => 
        \counter_points_snapshot[3]_net_1\, Y => 
        un4_data_in_validlt30_1);
    
    \counter_points_snapshot[13]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[13]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[13]_net_1\);
    
    \counter_points_snapshot[11]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[11]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[11]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I284_Y_0 : AX1A
      port map(A => N533, B => N529, C => 
        ADD_32x32_fast_I284_Y_0_0, Y => 
        \un1_data_out_valid_0_sqmuxa_2[4]\);
    
    \data_out[110]\ : DFN1C0
      port map(D => \sample_f0_wdata[46]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(110));
    
    \counter_points_snapshot_RNO_0[10]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[10]\, B => 
        nb_snapshot_param(10), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_96);
    
    \counter_points_snapshot_RNO[27]\ : XA1C
      port map(A => N746, B => ADD_32x32_fast_I307_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[27]\);
    
    \counter_points_snapshot[9]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[9]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[9]_net_1\);
    
    \counter_points_snapshot[28]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[28]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[28]_net_1\);
    
    \counter_points_snapshot_RNIVG9N[0]\ : NOR3C
      port map(A => un4_data_in_validlt30_2, B => 
        un4_data_in_validlt30_1, C => un4_data_in_validlt30_15, Y
         => un4_data_in_validlt30_23);
    
    \counter_points_snapshot_RNI37D9[24]\ : NOR2
      port map(A => \counter_points_snapshot[24]_net_1\, B => 
        \counter_points_snapshot[25]_net_1\, Y => 
        un4_data_in_validlt30_12);
    
    data_out_valid_0_sqmuxa : OR2B
      port map(A => sample_f0_val_0, B => start_snapshot_f0, Y
         => \data_out_valid_0_sqmuxa\);
    
    \counter_points_snapshot_RNO[19]\ : XA1B
      port map(A => N762, B => ADD_32x32_fast_I299_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[19]\);
    
    \data_out_RNO[96]\ : MX2
      port map(A => sample_f0_15, B => sample_f0_47, S => 
        data_shaping_R0_0, Y => \sample_f0_wdata[32]\);
    
    \data_out[91]\ : DFN1C0
      port map(D => \sample_f0_wdata[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(91));
    
    \data_out[120]\ : DFN1C0
      port map(D => sample_f0_wdata_56, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(120));
    
    \counter_points_snapshot_RNO[24]\ : XA1C
      port map(A => N752, B => ADD_32x32_fast_I304_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[24]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y : NOR3
      port map(A => N626, B => ADD_32x32_fast_I254_Y_0, C => N783, 
        Y => N746);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I190_Y : OR2
      port map(A => N586, B => N578, Y => N642);
    
    \data_out[130]\ : DFN1C0
      port map(D => sample_f0_wdata_66, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(130));
    
    \data_out[104]\ : DFN1C0
      port map(D => \sample_f0_wdata[40]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(104));
    
    \counter_points_snapshot_RNO_0[4]\ : MX2C
      port map(A => nb_snapshot_param(4), B => 
        \un1_data_out_valid_0_sqmuxa_2[4]\, S => 
        \counter_points_snapshot_2_sqmuxa\, Y => N_90);
    
    \counter_points_snapshot_RNIRK8P[14]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[14]_net_1\, Y => 
        \un1_counter_points_snapshot[17]\);
    
    \counter_points_snapshot_RNO_0[1]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[1]\, B => 
        nb_snapshot_param(1), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_87);
    
    \counter_points_snapshot_RNIHHQQ[3]\ : MX2
      port map(A => nb_snapshot_param(3), B => 
        \counter_points_snapshot[3]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[28]\);
    
    \data_out[102]\ : DFN1C0
      port map(D => \sample_f0_wdata[38]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(102));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I64_Y : AO1A
      port map(A => \un1_counter_points_snapshot[17]\, B => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, C => N419, Y => N507);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y : OR3B
      port map(A => ADD_32x32_fast_I252_Y_1, B => N777, C => N622, 
        Y => N742);
    
    \counter_points_snapshot_RNO[7]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_93, Y => 
        \counter_points_snapshot_10[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I309_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I309_Y_0_0);
    
    \counter_points_snapshot_RNO[12]\ : XA1B
      port map(A => N780, B => ADD_32x32_fast_I292_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[12]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I235_Y : OR2
      port map(A => N650, B => N634, Y => N771);
    
    \data_out[93]\ : DFN1C0
      port map(D => \sample_f0_wdata[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(93));
    
    \counter_points_snapshot_RNISO8P[15]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[15]_net_1\, Y => 
        \un1_counter_points_snapshot[16]\);
    
    \counter_points_snapshot[4]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[4]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[4]_net_1\);
    
    counter_points_snapshot_2_sqmuxa : OR3B
      port map(A => enable_f0, B => 
        \counter_points_snapshot_2_sqmuxa_2\, C => burst_f0, Y
         => \counter_points_snapshot_2_sqmuxa\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I301_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[10]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I301_Y_0_0);
    
    \data_out[159]\ : DFN1C0
      port map(D => sample_f0_wdata_95, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(159));
    
    \data_out[105]\ : DFN1C0
      port map(D => \sample_f0_wdata[41]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(105));
    
    \counter_points_snapshot[15]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[15]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[15]_net_1\);
    
    \data_out[141]\ : DFN1C0
      port map(D => sample_f0_wdata_77, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(141));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I108_Y : OR2
      port map(A => N495, B => N491, Y => N554);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I140_Y : OR2
      port map(A => N527, B => N523, Y => N586);
    
    \data_out[81]\ : DFN1C0
      port map(D => \sample_f0_wdata[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(81));
    
    \data_out_RNO[99]\ : MX2
      port map(A => sample_f0_12, B => sample_f0_44, S => 
        data_shaping_R0_0, Y => \sample_f0_wdata[35]\);
    
    \counter_points_snapshot_RNIB5QQ[0]\ : MX2
      port map(A => nb_snapshot_param(0), B => 
        \counter_points_snapshot[0]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1\, Y => 
        \un1_counter_points_snapshot[31]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I310_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I310_Y_0_0);
    
    \data_out_RNO[104]\ : MX2
      port map(A => sample_f0_7, B => sample_f0_39, S => 
        data_shaping_R0, Y => \sample_f0_wdata[40]\);
    
    \counter_points_snapshot[7]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[7]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[7]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y_0 : OR3
      port map(A => N487, B => N491, C => N558, Y => 
        ADD_32x32_fast_I256_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I234_Y_0_o2 : 
        NOR2
      port map(A => N771, B => I60_un1_Y, Y => N768);
    
    \data_out[114]\ : DFN1C0
      port map(D => sample_f0_wdata_50, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(114));
    
    \counter_points_snapshot_RNIR5RQ[8]\ : MX2C
      port map(A => nb_snapshot_param(8), B => 
        \counter_points_snapshot[8]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1\, Y => 
        \un1_counter_points_snapshot[23]\);
    
    \counter_points_snapshot[0]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[0]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[0]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I182_Y : OR3
      port map(A => N507, B => N511, C => N578, Y => N634);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I120_Y : OR2
      port map(A => N507, B => N503, Y => N566);
    
    \counter_points_snapshot[27]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[27]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[27]_net_1\);
    
    \data_out[143]\ : DFN1C0
      port map(D => sample_f0_wdata_79, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(143));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I199_Y : OR2
      port map(A => N590, B => N380, Y => N654);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I110_Y : OR2
      port map(A => ADD_32x32_fast_I110_Y_0, B => N497, Y => N556);
    
    \data_out[112]\ : DFN1C0
      port map(D => sample_f0_wdata_48, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(112));
    
    \counter_points_snapshot_RNIP88P[21]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[21]_net_1\, Y => 
        \un1_counter_points_snapshot[10]\);
    
    \data_out[124]\ : DFN1C0
      port map(D => sample_f0_wdata_60, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(124));
    
    \data_out[134]\ : DFN1C0
      port map(D => sample_f0_wdata_70, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(134));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I80_Y : OA1A
      port map(A => \un1_counter_points_snapshot[25]\, B => 
        \un1_counter_points_snapshot[26]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N523);
    
    \counter_points_snapshot_RNO[28]\ : XA1C
      port map(A => N744, B => ADD_32x32_fast_I308_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[28]\);
    
    \data_out[83]\ : DFN1C0
      port map(D => \sample_f0_wdata[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(83));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_2 : NOR3A
      port map(A => ADD_32x32_fast_I250_Y_1, B => N483, C => N487, 
        Y => ADD_32x32_fast_I250_Y_2);
    
    \data_out[122]\ : DFN1C0
      port map(D => sample_f0_wdata_58, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(122));
    
    \data_out[115]\ : DFN1C0
      port map(D => sample_f0_wdata_51, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(115));
    
    \counter_points_snapshot_RNID01S[10]\ : MX2C
      port map(A => nb_snapshot_param(10), B => 
        \counter_points_snapshot[10]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[21]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I44_Y : AOI1B
      port map(A => \un1_counter_points_snapshot[8]\, B => 
        \un1_counter_points_snapshot[7]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N487);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I38_Y_0_o2 : OA1
      port map(A => \un1_counter_points_snapshot[4]\, B => 
        \un1_counter_points_snapshot[5]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => I94_un1_Y);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y_0 : AOI1B
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        \un1_counter_points_snapshot[17]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I118_Y_0);
    
    \data_out[132]\ : DFN1C0
      port map(D => sample_f0_wdata_68, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(132));
    
    \counter_points_snapshot[30]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[30]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[30]_net_1\);
    
    \data_out[96]\ : DFN1C0
      port map(D => \sample_f0_wdata[32]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(96));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y : NOR3
      port map(A => N628, B => ADD_32x32_fast_I255_Y_0, C => N786, 
        Y => N748);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I294_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[17]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I294_Y_0_0);
    
    \data_out[125]\ : DFN1C0
      port map(D => sample_f0_wdata_61, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(125));
    
    \data_out[135]\ : DFN1C0
      port map(D => sample_f0_wdata_71, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(135));
    
    \data_out_RNO[87]\ : NOR2B
      port map(A => sample_f0_56, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[23]\);
    
    \data_out_RNO[108]\ : MX2
      port map(A => sample_f0_3, B => sample_f0_35, S => 
        data_shaping_R0, Y => \sample_f0_wdata[44]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I15_G0N : NOR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[16]\, Y => I60_un1_Y);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0 : NOR2
      port map(A => ADD_32x32_fast_I253_Y_0_0, B => N752, Y => 
        N744);
    
    \counter_points_snapshot_RNID9QQ[1]\ : MX2C
      port map(A => nb_snapshot_param(1), B => 
        \counter_points_snapshot[1]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1\, Y => 
        \un1_counter_points_snapshot[30]\);
    
    data_out_valid : DFN1C0
      port map(D => data_out_valid_19, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out_valid);
    
    \data_out_RNO[90]\ : NOR2B
      port map(A => sample_f0_53, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[26]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I174_Y : OR3
      port map(A => N507, B => N511, C => N562, Y => N626);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I29_G0N : OR3B
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1\, C => 
        data_out_valid_0_sqmuxa_1, Y => N467);
    
    \data_out[71]\ : DFN1C0
      port map(D => sample_f0_wdata_7, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(71));
    
    \data_out[65]\ : DFN1C0
      port map(D => sample_f0_wdata_1, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(65));
    
    \counter_points_snapshot_RNIUS8P[26]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[26]_net_1\, Y => 
        \un1_counter_points_snapshot[5]\);
    
    \counter_points_snapshot_RNIO88P[11]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[11]_net_1\, Y => 
        \un1_counter_points_snapshot[20]\);
    
    \counter_points_snapshot[18]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[18]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[18]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I260_Y : NOR3
      port map(A => N622, B => N638, C => N654, Y => N758);
    
    \data_out_RNO[98]\ : MX2
      port map(A => sample_f0_13, B => sample_f0_45, S => 
        data_shaping_R0_0, Y => \sample_f0_wdata[34]\);
    
    \data_out[86]\ : DFN1C0
      port map(D => \sample_f0_wdata[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(86));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I288_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[23]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I288_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I166_Y : OR2
      port map(A => N562, B => N554, Y => N618);
    
    \data_out[150]\ : DFN1C0
      port map(D => sample_f0_wdata_86, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(150));
    
    \counter_points_snapshot_RNIQC8P[22]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[22]_net_1\, Y => 
        \un1_counter_points_snapshot[9]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I297_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[17]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I297_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I296_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I296_Y_0_0);
    
    \data_out[148]\ : DFN1C0
      port map(D => sample_f0_wdata_84, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(148));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter_points_snapshot_RNIPC8P[12]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[12]_net_1\, Y => 
        \un1_counter_points_snapshot[19]\);
    
    \counter_points_snapshot_RNIB7E9[28]\ : NOR2
      port map(A => \counter_points_snapshot[28]_net_1\, B => 
        \counter_points_snapshot[29]_net_1\, Y => 
        un4_data_in_validlt30_14);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I13_G0N : NOR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[18]\, Y => N419);
    
    \counter_points_snapshot_RNIA0DC[6]\ : NOR3A
      port map(A => un4_data_in_validlt30_4, B => 
        \counter_points_snapshot[7]_net_1\, C => 
        \counter_points_snapshot[6]_net_1\, Y => 
        un4_data_in_validlt30_17);
    
    \counter_points_snapshot[8]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[8]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[8]_net_1\);
    
    counter_points_snapshot_2_sqmuxa_2 : NOR2A
      port map(A => start_snapshot_f0, B => sample_f0_val_0, Y
         => \counter_points_snapshot_2_sqmuxa_2\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I178_Y : OR2
      port map(A => N574, B => N566, Y => N630);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I136_Y : OR3
      port map(A => I74_un1_Y, B => N401, C => N523, Y => N582);
    
    \data_out[73]\ : DFN1C0
      port map(D => sample_f0_wdata_9, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(73));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I283_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[28]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I283_Y_0_0);
    
    \data_out[92]\ : DFN1C0
      port map(D => \sample_f0_wdata[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(92));
    
    \data_out[67]\ : DFN1C0
      port map(D => sample_f0_wdata_3, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(67));
    
    \data_out[107]\ : DFN1C0
      port map(D => \sample_f0_wdata[43]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(107));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y_0 : OR2
      port map(A => N644, B => N628, Y => ADD_32x32_fast_I263_Y_0);
    
    \counter_points_snapshot_RNO[6]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_92, Y => 
        \counter_points_snapshot_10[6]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I290_Y_0 : XNOR3
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[21]\, C => N786, Y => 
        \un1_data_out_valid_0_sqmuxa_2[10]\);
    
    \counter_points_snapshot[29]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[29]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[29]_net_1\);
    
    \counter_points_snapshot_RNIDBS75_1[31]\ : OR2B
      port map(A => data_out_valid_0_sqmuxa_1, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_data_out_valid_0_sqmuxa_1[31]\);
    
    \counter_points_snapshot_RNI28AJ4[31]\ : OR2
      port map(A => data_out_valid_0_sqmuxa_1_1, B => 
        un4_data_in_validlto30_i, Y => data_out_valid_0_sqmuxa_1);
    
    \data_out_RNO[94]\ : NOR2B
      port map(A => sample_f0_49, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[30]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I300_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[11]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I300_Y_0_0);
    
    \counter_points_snapshot_RNO[25]\ : XA1B
      port map(A => N750, B => ADD_32x32_fast_I305_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[25]\);
    
    \counter_points_snapshot[20]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[20]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[20]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I302_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[9]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I302_Y_0_0);
    
    \counter_points_snapshot_RNIR6C9[20]\ : NOR2
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        \counter_points_snapshot[21]_net_1\, Y => 
        un4_data_in_validlt30_10);
    
    \data_out_RNO[95]\ : NOR2B
      port map(A => sample_f0_48, B => data_shaping_R0, Y => 
        \sample_f0_wdata[31]\);
    
    \counter_points_snapshot[17]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[17]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[17]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I194_Y : OR2
      port map(A => N590, B => N582, Y => N646);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I88_Y : AOI1B
      port map(A => \un1_counter_points_snapshot[30]\, B => 
        \un1_counter_points_snapshot[29]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N531);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I292_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I292_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I28_G0N : OR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[3]\, Y => N464);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y : OR3A
      port map(A => ADD_32x32_fast_I250_Y_2, B => N618, C => N771, 
        Y => N738);
    
    \data_out_RNO[93]\ : NOR2B
      port map(A => sample_f0_50, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[29]\);
    
    \data_out[154]\ : DFN1C0
      port map(D => sample_f0_wdata_90, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(154));
    
    \counter_points_snapshot_RNITMC9[12]\ : NOR2
      port map(A => \counter_points_snapshot[12]_net_1\, B => 
        \counter_points_snapshot[13]_net_1\, Y => 
        un4_data_in_validlt30_6);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I261_Y_0_o2 : 
        OR2A
      port map(A => N764, B => N497, Y => N760);
    
    \data_out[82]\ : DFN1C0
      port map(D => \sample_f0_wdata[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(82));
    
    \data_out[117]\ : DFN1C0
      port map(D => sample_f0_wdata_53, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(117));
    
    \counter_points_snapshot_RNO[20]\ : XA1C
      port map(A => N760, B => ADD_32x32_fast_I300_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[20]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y_0 : OR3
      port map(A => N483, B => N487, C => N554, Y => 
        ADD_32x32_fast_I254_Y_0);
    
    \counter_points_snapshot_RNIT9RQ[9]\ : MX2C
      port map(A => nb_snapshot_param(9), B => 
        \counter_points_snapshot[9]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1\, Y => 
        \un1_counter_points_snapshot[22]\);
    
    \data_out[76]\ : DFN1C0
      port map(D => sample_f0_wdata_12, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(76));
    
    \data_out[152]\ : DFN1C0
      port map(D => sample_f0_wdata_88, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(152));
    
    \counter_points_snapshot_RNIVMC9[22]\ : NOR2
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        un4_data_in_validlt30_11);
    
    \data_out[149]\ : DFN1C0
      port map(D => sample_f0_wdata_85, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(149));
    
    \data_out[127]\ : DFN1C0
      port map(D => sample_f0_wdata_63, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(127));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I237_Y : NOR2
      port map(A => N654, B => N638, Y => N777);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I236_Y : OR2B
      port map(A => N652_i, B => N636, Y => N774);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I198_Y : NOR2
      port map(A => N588, B => N533, Y => N652_i);
    
    \data_out[137]\ : DFN1C0
      port map(D => sample_f0_wdata_73, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(137));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I30_G0N : OR3B
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => 
        data_out_valid_0_sqmuxa_1, Y => N470);
    
    \data_out_RNO[81]\ : NOR2B
      port map(A => sample_f0_62, B => data_shaping_R0, Y => 
        \sample_f0_wdata[17]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I144_Y : OR2
      port map(A => N531, B => N527, Y => N590);
    
    \data_out[155]\ : DFN1C0
      port map(D => sample_f0_wdata_91, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(155));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \counter_points_snapshot_RNO[5]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_91, Y => 
        \counter_points_snapshot_10[5]\);
    
    \counter_points_snapshot_RNO[17]\ : XA1B
      port map(A => N766, B => ADD_32x32_fast_I297_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[17]\);
    
    \counter_points_snapshot_RNI099P[19]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[19]_net_1\, Y => 
        \un1_counter_points_snapshot[12]\);
    
    data_out_valid_RNO_0 : AO1B
      port map(A => data_out_valid_0_sqmuxa_1, B => 
        \data_out_valid_0_sqmuxa\, C => enable_f0, Y => 
        un1_enable_2);
    
    \data_out[90]\ : DFN1C0
      port map(D => \sample_f0_wdata[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(90));
    
    \counter_points_snapshot[2]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[2]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[2]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y : OR3B
      port map(A => N620, B => ADD_32x32_fast_I251_Y_2, C => N774, 
        Y => N740);
    
    \counter_points_snapshot_RNO[14]\ : XA1C
      port map(A => N774, B => ADD_32x32_fast_I294_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[14]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I132_Y : OR3
      port map(A => I74_un1_Y, B => N401, C => N515, Y => N578);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I282_Y_0 : XNOR3
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[29]\, C => N533, Y => 
        \un1_data_out_valid_0_sqmuxa_2[2]\);
    
    \data_out_RNO[92]\ : NOR2B
      port map(A => sample_f0_51, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[28]\);
    
    \counter_points_snapshot_RNIO48P[20]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[20]_net_1\, Y => 
        \un1_counter_points_snapshot[11]\);
    
    \data_out[99]\ : DFN1C0
      port map(D => \sample_f0_wdata[35]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(99));
    
    \data_out_RNO[100]\ : MX2
      port map(A => sample_f0_11, B => sample_f0_43, S => 
        data_shaping_R0, Y => \sample_f0_wdata[36]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I258_Y : NOR3
      port map(A => N634, B => N618, C => N650, Y => N754);
    
    \counter_points_snapshot_RNISK8P[24]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[24]_net_1\, Y => 
        \un1_counter_points_snapshot[7]\);
    
    \data_out[106]\ : DFN1C0
      port map(D => \sample_f0_wdata[42]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(106));
    
    \counter_points_snapshot_RNO[21]\ : XA1C
      port map(A => N758, B => ADD_32x32_fast_I301_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[21]\);
    
    \counter_points_snapshot_RNITO8P[25]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[25]_net_1\, Y => 
        \un1_counter_points_snapshot[6]\);
    
    \counter_points_snapshot_RNITNQ14[6]\ : NOR3C
      port map(A => un4_data_in_validlt30_26, B => 
        un4_data_in_validlt30_25, C => un4_data_in_validlt30_27, 
        Y => un4_data_in_validlto30_i);
    
    \data_out_RNO[103]\ : MX2
      port map(A => sample_f0_8, B => sample_f0_40, S => 
        data_shaping_R0, Y => \sample_f0_wdata[39]\);
    
    \counter_points_snapshot_RNIVEFM1[6]\ : NOR3C
      port map(A => un4_data_in_validlt30_18, B => 
        un4_data_in_validlt30_17, C => un4_data_in_validlt30_23, 
        Y => un4_data_in_validlt30_27);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I128_Y : OR2
      port map(A => N515, B => N511, Y => N574);
    
    \data_out[98]\ : DFN1C0
      port map(D => \sample_f0_wdata[34]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(98));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y : NOR3
      port map(A => I60_un1_Y, B => N431, C => 
        ADD_32x32_fast_I118_Y_0, Y => N564);
    
    \counter_points_snapshot_RNIFDQQ[2]\ : MX2C
      port map(A => nb_snapshot_param(2), B => 
        \counter_points_snapshot[2]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[29]\);
    
    \data_out[80]\ : DFN1C0
      port map(D => \sample_f0_wdata[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(80));
    
    \data_out[72]\ : DFN1C0
      port map(D => sample_f0_wdata_8, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(72));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y : NOR3
      port map(A => N630, B => ADD_32x32_fast_I256_Y_0, C => N789, 
        Y => N750);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I288_Y_0 : AX1B
      port map(A => N401, B => N650, C => 
        ADD_32x32_fast_I288_Y_0_0, Y => 
        \un1_data_out_valid_0_sqmuxa_2[8]\);
    
    \data_out_RNO[107]\ : MX2
      port map(A => sample_f0_4, B => sample_f0_36, S => 
        data_shaping_R0, Y => \sample_f0_wdata[43]\);
    
    \data_out[89]\ : DFN1C0
      port map(D => \sample_f0_wdata[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(89));
    
    \counter_points_snapshot_RNI059P[28]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[28]_net_1\, Y => 
        \un1_counter_points_snapshot[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y : NOR2
      port map(A => ADD_32x32_fast_I263_Y_0, B => N533, Y => N764);
    
    \counter_points_snapshot_RNIQG8P[13]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[13]_net_1\, Y => 
        \un1_counter_points_snapshot[18]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I289_Y_0 : XNOR2
      port map(A => ADD_32x32_fast_I289_Y_0_0, B => N789, Y => 
        \un1_data_out_valid_0_sqmuxa_2[9]\);
    
    \data_out_RNO[101]\ : MX2
      port map(A => sample_f0_10, B => sample_f0_42, S => 
        data_shaping_R0, Y => \sample_f0_wdata[37]\);
    
    \data_out[116]\ : DFN1C0
      port map(D => sample_f0_wdata_52, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(116));
    
    \counter_points_snapshot[19]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[19]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[19]_net_1\);
    
    \counter_points_snapshot_RNO_0[2]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[2]\, B => 
        nb_snapshot_param(2), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_88);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I298_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[13]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I298_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I197_Y : OR2
      port map(A => N594, B => N586, Y => N650);
    
    \counter_points_snapshot_RNITS8P[16]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1\, B => 
        \counter_points_snapshot[16]_net_1\, Y => 
        \un1_counter_points_snapshot[15]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I285_Y_0 : XOR3
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[26]\, C => N654, Y => 
        \un1_data_out_valid_0_sqmuxa_2[5]\);
    
    \counter_points_snapshot[10]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[10]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[10]_net_1\);
    
    \counter_points_snapshot_RNO[18]\ : XA1C
      port map(A => N764, B => ADD_32x32_fast_I298_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[18]\);
    
    \data_out[88]\ : DFN1C0
      port map(D => \sample_f0_wdata[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(88));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_S_0 : XOR2
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[31]\, Y => 
        \un1_data_out_valid_0_sqmuxa_2[0]\);
    
    \data_out[126]\ : DFN1C0
      port map(D => sample_f0_wdata_62, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(126));
    
    \data_out[94]\ : DFN1C0
      port map(D => \sample_f0_wdata[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(94));
    
    \data_out[140]\ : DFN1C0
      port map(D => sample_f0_wdata_76, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(140));
    
    \data_out[136]\ : DFN1C0
      port map(D => sample_f0_wdata_72, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(136));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I27_G0N : OR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[4]\, Y => N461);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I293_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[18]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I293_Y_0_0);
    
    \counter_points_snapshot[22]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[22]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[22]_net_1\);
    
    \data_out_RNO[86]\ : NOR2B
      port map(A => sample_f0_57, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[22]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I147_Y : OR2
      port map(A => N531, B => N380, Y => N594);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I304_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[7]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I304_Y_0_0);
    
    data_out_valid_RNO_1 : NOR2B
      port map(A => enable_f0, B => burst_f0, Y => 
        counter_points_snapshot_0_sqmuxa_i);
    
    \data_out[101]\ : DFN1C0
      port map(D => \sample_f0_wdata[37]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(101));
    
    \data_out[157]\ : DFN1C0
      port map(D => sample_f0_wdata_93, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(157));
    
    \counter_points_snapshot_RNO[4]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_90, Y => 
        \counter_points_snapshot_10[4]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I110_Y_0 : OA1A
      port map(A => \un1_counter_points_snapshot[11]\, B => 
        \un1_counter_points_snapshot[10]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I110_Y_0);
    
    \counter_points_snapshot_RNO[30]\ : XA1B
      port map(A => N740, B => ADD_32x32_fast_I310_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[30]\);
    
    \counter_points_snapshot[6]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[6]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[6]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I54_Y_0_o2 : 
        AO1C
      port map(A => \un1_counter_points_snapshot[12]\, B => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, C => N434, Y => N497);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I176_Y : OR2A
      port map(A => N564, B => N572, Y => N628);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y_0 : AO1B
      port map(A => \un1_counter_points_snapshot[25]\, B => 
        \un1_counter_points_snapshot[23]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I134_Y_0);
    
    \data_out[70]\ : DFN1C0
      port map(D => sample_f0_wdata_6, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(70));
    
    \counter_points_snapshot_RNO_0[5]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[5]\, B => 
        nb_snapshot_param(5), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_91);
    
    \data_out[84]\ : DFN1C0
      port map(D => \sample_f0_wdata[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(84));
    
    \data_out[103]\ : DFN1C0
      port map(D => \sample_f0_wdata[39]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(103));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I7_G0N : NOR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[24]\, Y => N401);
    
    \counter_points_snapshot_RNIRG8P[23]\ : OR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        \un1_counter_points_snapshot[8]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I84_Y : OA1
      port map(A => \un1_counter_points_snapshot[28]\, B => 
        \un1_counter_points_snapshot[27]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N527);
    
    \counter_points_snapshot[5]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[5]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[5]_net_1\);
    
    \counter_points_snapshot_RNO[26]\ : XA1C
      port map(A => N748, B => ADD_32x32_fast_I306_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[26]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I8_G0N : NOR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[23]\, Y => I74_un1_Y);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I289_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[22]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I289_Y_0_0);
    
    \data_out[79]\ : DFN1C0
      port map(D => sample_f0_wdata_15, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(79));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I281_Y_0 : XNOR3
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[30]\, C => N380, Y => 
        \un1_data_out_valid_0_sqmuxa_2[1]\);
    
    \data_out[144]\ : DFN1C0
      port map(D => sample_f0_wdata_80, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(144));
    
    \data_out_RNO[89]\ : NOR2B
      port map(A => sample_f0_54, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[25]\);
    
    \counter_points_snapshot_RNO[8]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_94, Y => 
        \counter_points_snapshot_10[8]\);
    
    \data_out[111]\ : DFN1C0
      port map(D => \sample_f0_wdata[47]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(111));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I295_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[16]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I295_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_CO1 : NOR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[31]\, Y => N380);
    
    \data_out[142]\ : DFN1C0
      port map(D => sample_f0_wdata_78, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(142));
    
    \data_out[78]\ : DFN1C0
      port map(D => sample_f0_wdata_14, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(78));
    
    \counter_points_snapshot_RNO[23]\ : XA1B
      port map(A => N754, B => ADD_32x32_fast_I303_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[23]\);
    
    \counter_points_snapshot_RNIDBS75[31]\ : OR2B
      port map(A => data_out_valid_0_sqmuxa_1, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I184_Y : NOR2
      port map(A => N580, B => N572, Y => N636);
    
    \counter_points_snapshot_RNO_0[3]\ : MX2C
      port map(A => nb_snapshot_param(3), B => 
        \un1_data_out_valid_0_sqmuxa_2[3]\, S => 
        \counter_points_snapshot_2_sqmuxa\, Y => N_89);
    
    \counter_points_snapshot_RNI5HSA[0]\ : NOR3
      port map(A => \counter_points_snapshot[1]_net_1\, B => 
        \counter_points_snapshot[0]_net_1\, C => 
        \counter_points_snapshot[30]_net_1\, Y => 
        un4_data_in_validlt30_15);
    
    \counter_points_snapshot[26]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[26]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[26]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I305_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[6]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I305_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y_1 : NOR3A
      port map(A => ADD_32x32_fast_I252_Y_0, B => N487, C => N491, 
        Y => ADD_32x32_fast_I252_Y_1);
    
    \data_out[121]\ : DFN1C0
      port map(D => sample_f0_wdata_57, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(121));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I60_Y : AO1A
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, C => I60_un1_Y, Y
         => N503);
    
    \counter_points_snapshot_RNO[0]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_86, Y => 
        \counter_points_snapshot_10[0]\);
    
    \data_out[131]\ : DFN1C0
      port map(D => sample_f0_wdata_67, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(131));
    
    \data_out[113]\ : DFN1C0
      port map(D => sample_f0_wdata_49, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(113));
    
    \data_out[145]\ : DFN1C0
      port map(D => sample_f0_wdata_81, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(145));
    
    \counter_points_snapshot_RNI5ND9[16]\ : NOR2
      port map(A => \counter_points_snapshot[16]_net_1\, B => 
        \counter_points_snapshot[17]_net_1\, Y => 
        un4_data_in_validlt30_8);
    
    \counter_points_snapshot_RNIIURI[26]\ : NOR3A
      port map(A => un4_data_in_validlt30_14, B => 
        \counter_points_snapshot[27]_net_1\, C => 
        \counter_points_snapshot[26]_net_1\, Y => 
        un4_data_in_validlt30_22);
    
    \data_out[66]\ : DFN1C0
      port map(D => sample_f0_wdata_2, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(66));
    
    \counter_points_snapshot[1]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[1]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[1]_net_1\);
    
    \counter_points_snapshot_RNO[31]\ : XA1C
      port map(A => N738, B => ADD_32x32_fast_I311_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[31]\);
    
    \data_out_RNO[109]\ : MX2
      port map(A => sample_f0_2, B => sample_f0_34, S => 
        data_shaping_R0, Y => \sample_f0_wdata[45]\);
    
    \counter_points_snapshot_RNO_0[0]\ : MX2C
      port map(A => nb_snapshot_param(0), B => 
        \un1_data_out_valid_0_sqmuxa_2[0]\, S => 
        \counter_points_snapshot_2_sqmuxa\, Y => N_86);
    
    \counter_points_snapshot_RNO[15]\ : XA1C
      port map(A => N771, B => ADD_32x32_fast_I295_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[15]\);
    
    \data_out[123]\ : DFN1C0
      port map(D => sample_f0_wdata_59, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(123));
    
    \counter_points_snapshot_RNIKSL51[22]\ : NOR3C
      port map(A => un4_data_in_validlt30_12, B => 
        un4_data_in_validlt30_11, C => un4_data_in_validlt30_22, 
        Y => un4_data_in_validlt30_26);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    counter_points_snapshot_3_sqmuxa : OR2
      port map(A => start_snapshot_f0, B => burst_f0, Y => 
        \counter_points_snapshot_3_sqmuxa\);
    
    \data_out[133]\ : DFN1C0
      port map(D => sample_f0_wdata_69, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(133));
    
    \counter_points_snapshot_RNIACL51[14]\ : NOR3C
      port map(A => un4_data_in_validlt30_8, B => 
        un4_data_in_validlt30_7, C => un4_data_in_validlt30_20, Y
         => un4_data_in_validlt30_25);
    
    \counter_points_snapshot_RNO[29]\ : XA1B
      port map(A => N742, B => ADD_32x32_fast_I309_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[29]\);
    
    \counter_points_snapshot_RNIVF66[4]\ : NOR2
      port map(A => \counter_points_snapshot[4]_net_1\, B => 
        \counter_points_snapshot[5]_net_1\, Y => 
        un4_data_in_validlt30_2);
    
    \counter_points_snapshot[31]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[31]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[31]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I36_Y : OR2B
      port map(A => N464, B => N461, Y => N479);
    
    \data_out_RNO[97]\ : MX2
      port map(A => sample_f0_14, B => sample_f0_46, S => 
        data_shaping_R0_0, Y => \sample_f0_wdata[33]\);
    
    \data_out[74]\ : DFN1C0
      port map(D => sample_f0_wdata_10, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(74));
    
    \counter_points_snapshot_RNO[10]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_96, Y => 
        \counter_points_snapshot_10[10]\);
    
    \data_out[108]\ : DFN1C0
      port map(D => \sample_f0_wdata[44]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(108));
    
    \counter_points_snapshot_RNO_0[6]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[6]\, B => 
        nb_snapshot_param(6), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_92);
    
    \data_out[156]\ : DFN1C0
      port map(D => sample_f0_wdata_92, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(156));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I240_Y : OR2
      port map(A => N644, B => N533, Y => N786);
    
    \data_out_RNO[106]\ : MX2
      port map(A => sample_f0_5, B => sample_f0_37, S => 
        data_shaping_R0, Y => \sample_f0_wdata[42]\);
    
    \counter_points_snapshot_RNO_0[8]\ : MX2C
      port map(A => \un1_data_out_valid_0_sqmuxa_2[8]\, B => 
        nb_snapshot_param(8), S => 
        \counter_points_snapshot_2_sqmuxa_2\, Y => N_94);
    
    \data_out_RNO[80]\ : NOR2B
      port map(A => sample_f0_63, B => data_shaping_R0, Y => 
        \sample_f0_wdata[16]\);
    
    \counter_points_snapshot_RNO[1]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_87, Y => 
        \counter_points_snapshot_10[1]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I303_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[8]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I303_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I40_Y : OA1A
      port map(A => \un1_counter_points_snapshot[6]\, B => 
        \un1_counter_points_snapshot[5]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N483);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I257_Y_0_o2 : 
        OR2
      port map(A => N756, B => N489, Y => N752);
    
    \counter_points_snapshot_RNO[22]\ : XA1C
      port map(A => N756, B => ADD_32x32_fast_I302_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[22]\);
    
    \data_out_RNO[88]\ : NOR2B
      port map(A => sample_f0_55, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[24]\);
    
    \counter_points_snapshot[12]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[12]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[12]_net_1\);
    
    \counter_points_snapshot[24]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[24]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[24]_net_1\);
    
    \data_out[95]\ : DFN1C0
      port map(D => \sample_f0_wdata[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(95));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y_0 : NOR2
      port map(A => N479, B => N483, Y => ADD_32x32_fast_I252_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y : OR3A
      port map(A => ADD_32x32_fast_I126_Y_1, B => N419, C => 
        I66_un1_Y, Y => N572);
    
    \data_out_RNO[110]\ : MX2
      port map(A => sample_f0_1, B => sample_f0_33, S => 
        data_shaping_R0, Y => \sample_f0_wdata[46]\);
    
    \counter_points_snapshot_RNO_0[9]\ : MX2C
      port map(A => nb_snapshot_param(9), B => 
        \un1_data_out_valid_0_sqmuxa_2[9]\, S => 
        \counter_points_snapshot_2_sqmuxa\, Y => N_95);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y_1 : AO1C
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        \un1_counter_points_snapshot[21]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I126_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I116_Y : OR3A
      port map(A => N434, B => N431, C => N503, Y => N562);
    
    \counter_points_snapshot_RNO[3]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_89, Y => 
        \counter_points_snapshot_10[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y_0 : OAI1
      port map(A => \un1_counter_points_snapshot[27]\, B => 
        \un1_counter_points_snapshot[26]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I142_Y_0);
    
    \data_out[118]\ : DFN1C0
      port map(D => sample_f0_wdata_54, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(118));
    
    counter_points_snapshot_0_sqmuxa_1_0 : OR2
      port map(A => \data_out_valid_0_sqmuxa\, B => burst_f0, Y
         => \counter_points_snapshot_0_sqmuxa_1_0\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I241_Y : OR2
      port map(A => N646, B => N380, Y => N789);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I306_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[5]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I306_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_1 : NOR3B
      port map(A => N467, B => N464, C => I94_un1_Y, Y => 
        ADD_32x32_fast_I251_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I239_Y : OR2
      port map(A => N642, B => N594, Y => N783);
    
    \counter_points_snapshot_RNIDBS75_0[31]\ : OR2B
      port map(A => data_out_valid_0_sqmuxa_1, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I287_Y_0 : XOR2
      port map(A => ADD_32x32_fast_I287_Y_0_0, B => N650, Y => 
        \un1_data_out_valid_0_sqmuxa_2[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I286_Y_0 : XOR3
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[25]\, C => N652_i, Y => 
        \un1_data_out_valid_0_sqmuxa_2[6]\);
    
    \counter_points_snapshot_RNIV09P[27]\ : NOR2B
      port map(A => \counter_points_snapshot_0_sqmuxa_1_0\, B => 
        \counter_points_snapshot[27]_net_1\, Y => 
        \un1_counter_points_snapshot[4]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I46_Y_0_o2 : 
        AOI1B
      port map(A => \un1_counter_points_snapshot[8]\, B => 
        \un1_counter_points_snapshot[9]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => N489);
    
    \data_out[128]\ : DFN1C0
      port map(D => sample_f0_wdata_64, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(128));
    
    \counter_points_snapshot_RNO[11]\ : XA1B
      port map(A => N783, B => ADD_32x32_fast_I291_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[11]\);
    
    \data_out[97]\ : DFN1C0
      port map(D => \sample_f0_wdata[33]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(97));
    
    \data_out[138]\ : DFN1C0
      port map(D => sample_f0_wdata_74, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(138));
    
    \data_out_RNO[84]\ : NOR2B
      port map(A => sample_f0_59, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[20]\);
    
    \data_out[85]\ : DFN1C0
      port map(D => \sample_f0_wdata[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(85));
    
    \counter_points_snapshot[3]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[3]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[3]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I18_G0N : OR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[13]\, Y => N434);
    
    \data_out_RNO[85]\ : NOR2B
      port map(A => sample_f0_58, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[21]\);
    
    \data_out[109]\ : DFN1C0
      port map(D => \sample_f0_wdata[45]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(109));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I259_Y_0 : NOR2B
      port map(A => N636, B => N620, Y => ADD_32x32_fast_I259_Y_0);
    
    \counter_points_snapshot_RNI4EQI[18]\ : NOR3A
      port map(A => un4_data_in_validlt30_10, B => 
        \counter_points_snapshot[19]_net_1\, C => 
        \counter_points_snapshot[18]_net_1\, Y => 
        un4_data_in_validlt30_20);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I68_Y : AO1
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[20]\, C => I66_un1_Y, Y => 
        N511);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I192_Y : OR2
      port map(A => N588, B => N580, Y => N644);
    
    \data_out_RNO[111]\ : MX2
      port map(A => sample_f0_0, B => sample_f0_32, S => 
        data_shaping_R0, Y => \sample_f0_wdata[47]\);
    
    \counter_points_snapshot[23]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[23]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[23]_net_1\);
    
    \counter_points_snapshot[21]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[21]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[21]_net_1\);
    
    \counter_points_snapshot[16]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[16]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[16]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y_0 : OR3
      port map(A => N485, B => N489, C => N556, Y => 
        ADD_32x32_fast_I255_Y_0);
    
    \data_out[147]\ : DFN1C0
      port map(D => sample_f0_wdata_83, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(147));
    
    \data_out[151]\ : DFN1C0
      port map(D => sample_f0_wdata_87, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(151));
    
    \data_out_RNO[83]\ : NOR2B
      port map(A => sample_f0_60, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[19]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I299_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[12]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I299_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I308_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[3]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I308_Y_0_0);
    
    \data_out[87]\ : DFN1C0
      port map(D => \sample_f0_wdata[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(87));
    
    \data_out[153]\ : DFN1C0
      port map(D => sample_f0_wdata_89, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(153));
    
    \counter_points_snapshot_RNIP1RQ[7]\ : MX2
      port map(A => nb_snapshot_param(7), B => 
        \counter_points_snapshot[7]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1\, Y => 
        \un1_counter_points_snapshot[24]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I283_Y_0 : XOR2
      port map(A => ADD_32x32_fast_I283_Y_0_0, B => N594, Y => 
        \un1_data_out_valid_0_sqmuxa_2[3]\);
    
    \counter_points_snapshot_RNI17D9[14]\ : NOR2
      port map(A => \counter_points_snapshot[14]_net_1\, B => 
        \counter_points_snapshot[15]_net_1\, Y => 
        un4_data_in_validlt30_7);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I259_Y : OR2B
      port map(A => ADD_32x32_fast_I259_Y_0, B => N652_i, Y => 
        N756);
    
    counter_points_snapshot_0_sqmuxa_1 : OR2
      port map(A => \data_out_valid_0_sqmuxa\, B => burst_f0, Y
         => \counter_points_snapshot_0_sqmuxa_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I86_Y : AO1C
      port map(A => \un1_counter_points_snapshot[28]\, B => 
        \un1_counter_points_snapshot[29]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N529);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y : OR2B
      port map(A => ADD_32x32_fast_I142_Y_0, B => N529, Y => N588);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I307_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[4]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I307_Y_0_0);
    
    \data_out_RNO[91]\ : NOR2B
      port map(A => sample_f0_52, B => data_shaping_R0_0, Y => 
        \sample_f0_wdata[27]\);
    
    \data_out[119]\ : DFN1C0
      port map(D => sample_f0_wdata_55, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(119));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_1 : NOR3B
      port map(A => N467, B => N470, C => N479, Y => 
        ADD_32x32_fast_I250_Y_1);
    
    \data_out_RNO[102]\ : MX2
      port map(A => sample_f0_9, B => sample_f0_41, S => 
        data_shaping_R0, Y => \sample_f0_wdata[38]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I72_Y : AO1A
      port map(A => \un1_counter_points_snapshot[21]\, B => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, C => N407, Y => N515);
    
    \counter_points_snapshot_RNILPQQ[5]\ : MX2
      port map(A => nb_snapshot_param(5), B => 
        \counter_points_snapshot[5]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[26]\);
    
    \counter_points_snapshot_RNO_0[7]\ : MX2C
      port map(A => nb_snapshot_param(7), B => 
        \un1_data_out_valid_0_sqmuxa_2[7]\, S => 
        \counter_points_snapshot_2_sqmuxa\, Y => N_93);
    
    \counter_points_snapshot_RNO[9]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_95, Y => 
        \counter_points_snapshot_10[9]\);
    
    \counter_points_snapshot_RNI5GFH[31]\ : OR3A
      port map(A => sample_f0_val_0, B => start_snapshot_f0, C
         => \counter_points_snapshot[31]_net_1\, Y => 
        data_out_valid_0_sqmuxa_1_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I291_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I291_Y_0_0);
    
    \data_out[69]\ : DFN1C0
      port map(D => sample_f0_wdata_5, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(69));
    
    \data_out[129]\ : DFN1C0
      port map(D => sample_f0_wdata_65, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(129));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I112_Y : OR3A
      port map(A => N434, B => N431, C => N495, Y => N558);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I311_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[31]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I311_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_2 : NOR3A
      port map(A => ADD_32x32_fast_I251_Y_1, B => N485, C => N489, 
        Y => ADD_32x32_fast_I251_Y_2);
    
    \data_out[139]\ : DFN1C0
      port map(D => sample_f0_wdata_75, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(139));
    
    \counter_points_snapshot[25]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[25]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[25]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I48_Y : OA1A
      port map(A => \un1_counter_points_snapshot[9]\, B => 
        \un1_counter_points_snapshot[10]\, C => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => N491);
    
    \data_out_RNO[82]\ : NOR2B
      port map(A => sample_f0_61, B => data_shaping_R0, Y => 
        \sample_f0_wdata[18]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y : OR3A
      port map(A => ADD_32x32_fast_I134_Y_0, B => N401, C => N407, 
        Y => N580);
    
    \counter_points_snapshot_RNIMTOI[10]\ : NOR3A
      port map(A => un4_data_in_validlt30_6, B => 
        \counter_points_snapshot[11]_net_1\, C => 
        \counter_points_snapshot[10]_net_1\, Y => 
        un4_data_in_validlt30_18);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I238_Y_0_o2 : 
        AO1
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[20]\, C => N783, Y => N780);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I90_Y : AO1A
      port map(A => \un1_counter_points_snapshot[30]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, C => N380, Y => 
        N533);
    
    \counter_points_snapshot_RNIJLQQ[4]\ : MX2
      port map(A => nb_snapshot_param(4), B => 
        \counter_points_snapshot[4]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[27]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I42_Y : AOI1B
      port map(A => \un1_counter_points_snapshot[7]\, B => 
        \un1_counter_points_snapshot[6]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N485);
    
    \counter_points_snapshot_RNI7G66[8]\ : NOR2
      port map(A => \counter_points_snapshot[8]_net_1\, B => 
        \counter_points_snapshot[9]_net_1\, Y => 
        un4_data_in_validlt30_4);
    
    un1_counter_points_snapshot_0_sqmuxa_1 : AO1B
      port map(A => \counter_points_snapshot_3_sqmuxa\, B => 
        \counter_points_snapshot_0_sqmuxa_1_0\, C => enable_f0, Y
         => un1_counter_points_snapshot_0_sqmuxa_1_i);
    
    \data_out[75]\ : DFN1C0
      port map(D => sample_f0_wdata_11, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(75));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I284_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[27]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_1[31]\, Y => 
        ADD_32x32_fast_I284_Y_0_0);
    
    \data_out[68]\ : DFN1C0
      port map(D => sample_f0_wdata_4, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(68));
    
    \counter_points_snapshot[14]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[14]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[14]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I12_G0N : NOR2B
      port map(A => \un1_data_out_valid_0_sqmuxa_1[31]\, B => 
        \un1_counter_points_snapshot[19]\, Y => I66_un1_Y);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I52_Y : AOI1B
      port map(A => \un1_counter_points_snapshot[12]\, B => 
        \un1_counter_points_snapshot[11]\, C => 
        \un1_data_out_valid_0_sqmuxa_1[31]\, Y => N495);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I168_Y : NOR2A
      port map(A => N564, B => N556, Y => N620);
    
    \counter_points_snapshot_RNINTQQ[6]\ : MX2C
      port map(A => nb_snapshot_param(6), B => 
        \counter_points_snapshot[6]_net_1\, S => 
        \counter_points_snapshot_0_sqmuxa_1_0\, Y => 
        \un1_counter_points_snapshot[25]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I264_Y : NOR3
      port map(A => N646, B => N380, C => N630, Y => N766);
    
    \counter_points_snapshot_RNO[16]\ : XA1B
      port map(A => N768, B => ADD_32x32_fast_I296_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[16]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I170_Y : OR2
      port map(A => N566, B => N558, Y => N622);
    
    data_out_valid_RNO : MX2A
      port map(A => un1_enable_2, B => sample_f0_val_0, S => 
        counter_points_snapshot_0_sqmuxa_i, Y => 
        data_out_valid_19);
    
    \data_out[100]\ : DFN1C0
      port map(D => \sample_f0_wdata[36]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(100));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I9_G0N : NOR2A
      port map(A => \un1_data_out_valid_0_sqmuxa_1_1[31]\, B => 
        \un1_counter_points_snapshot[22]\, Y => N407);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I262_Y : NOR3
      port map(A => N642, B => N594, C => N626, Y => N762);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0_0 : OR2
      port map(A => I94_un1_Y, B => N485, Y => 
        ADD_32x32_fast_I253_Y_0_0);
    
    \data_out[77]\ : DFN1C0
      port map(D => sample_f0_wdata_13, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(77));
    
    \data_out[146]\ : DFN1C0
      port map(D => sample_f0_wdata_82, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(146));
    
    \counter_points_snapshot_RNO[2]\ : NOR3A
      port map(A => enable_f0, B => burst_f0, C => N_88, Y => 
        \counter_points_snapshot_10[2]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I186_Y : OR2
      port map(A => N582, B => N574, Y => N638);
    
    \counter_points_snapshot_RNO[13]\ : XA1C
      port map(A => N777, B => ADD_32x32_fast_I293_Y_0_0, C => 
        un1_counter_points_snapshot_0_sqmuxa_1_i, Y => 
        \counter_points_snapshot_10[13]\);
    
    \data_out[158]\ : DFN1C0
      port map(D => sample_f0_wdata_94, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(158));
    
    \data_out_RNO[105]\ : MX2
      port map(A => sample_f0_6, B => sample_f0_38, S => 
        data_shaping_R0, Y => \sample_f0_wdata[41]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I17_G0N : NOR3B
      port map(A => \counter_points_snapshot[17]_net_1\, B => 
        \counter_points_snapshot_0_sqmuxa_1\, C => 
        data_out_valid_0_sqmuxa_1, Y => N431);
    
    \data_out[64]\ : DFN1C0
      port map(D => sample_f0_wdata_0, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f0_out(64));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I287_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[24]\, B => 
        \un1_data_out_valid_0_sqmuxa_1_0[31]\, Y => 
        ADD_32x32_fast_I287_Y_0_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1 is

    port( sample_f2_wdata   : in    std_logic_vector(95 downto 0);
          data_f2_out       : out   std_logic_vector(159 downto 64);
          nb_snapshot_param : in    std_logic_vector(0 to 0);
          HRESETn_c         : in    std_logic;
          HCLK_c            : in    std_logic;
          data_f2_out_valid : out   std_logic;
          I_13_20           : in    std_logic;
          I_9_20            : in    std_logic;
          I_5_20            : in    std_logic;
          I_38_4            : in    std_logic;
          I_31_5            : in    std_logic;
          N_4               : in    std_logic;
          I_45_4            : in    std_logic;
          I_56_4            : in    std_logic;
          I_52_4            : in    std_logic;
          I_24_4            : in    std_logic;
          I_20_12           : in    std_logic;
          enable_f2         : in    std_logic;
          burst_f2          : in    std_logic;
          start_snapshot_f2 : in    std_logic;
          sample_f2_val     : in    std_logic
        );

end lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1;

architecture DEF_ARCH of 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal counter_points_snapshot_0_sqmuxa_1_0, N_47_1, 
        un1_data_in_valid, 
        \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, N_47_0, 
        ADD_32x32_fast_I311_Y_0_0, 
        \counter_points_snapshot[31]_net_1\, 
        ADD_32x32_fast_I296_Y_0_0, 
        \un1_counter_points_snapshot[15]\, 
        ADD_32x32_fast_I250_Y_3, ADD_32x32_fast_I250_Y_1, N618, 
        N546, I32_un1_Y, N470, N479, ADD_32x32_fast_I308_Y_0_0, 
        \un1_counter_points_snapshot[3]\, 
        ADD_32x32_fast_I295_Y_0_0, 
        \counter_points_snapshot[15]_net_1\, 
        ADD_32x32_fast_I310_Y_0_0, 
        \counter_points_snapshot[30]_net_1\, 
        ADD_32x32_fast_I303_Y_0_0, 
        \un1_counter_points_snapshot[8]\, 
        ADD_32x32_fast_I304_Y_0_0, 
        \un1_counter_points_snapshot[7]\, 
        ADD_32x32_fast_I253_Y_0_0, N461, N458, N485, 
        ADD_32x32_fast_I307_Y_0_0, 
        \counter_points_snapshot[27]_net_1\, 
        ADD_32x32_fast_I292_Y_0_0, 
        \un1_counter_points_snapshot[19]\, 
        ADD_32x32_fast_I309_Y_0_0, 
        \counter_points_snapshot[29]_net_1\, 
        ADD_32x32_fast_I300_Y_0_0, 
        \counter_points_snapshot[20]_net_1\, 
        ADD_32x32_fast_I287_Y_0_0, 
        \un1_counter_points_snapshot[24]\, 
        ADD_32x32_fast_I251_Y_2, ADD_32x32_fast_I251_Y_1, N489, 
        ADD_32x32_fast_I251_Y_0, ADD_32x32_fast_I305_Y_0_0, 
        \counter_points_snapshot[25]_net_1\, 
        ADD_32x32_fast_I302_Y_0_0, 
        \counter_points_snapshot[22]_net_1\, 
        ADD_32x32_fast_I294_Y_0_0, 
        \un1_counter_points_snapshot[17]\, 
        ADD_32x32_fast_I299_Y_0_0, 
        \un1_counter_points_snapshot[12]\, 
        ADD_32x32_fast_I306_Y_0_0, 
        \counter_points_snapshot[26]_net_1\, 
        ADD_32x32_fast_I254_Y_0, N554, ADD_32x32_fast_I301_Y_0_0, 
        \counter_points_snapshot[21]_net_1\, 
        ADD_32x32_fast_I297_Y_0_0, 
        \un1_counter_points_snapshot[14]\, 
        ADD_32x32_fast_I252_Y_1, N483, N550, 
        ADD_32x32_fast_I298_Y_0_0, 
        \un1_counter_points_snapshot[13]\, 
        ADD_32x32_fast_I293_Y_0_0, 
        \counter_points_snapshot[13]_net_1\, 
        ADD_32x32_fast_I256_Y_0, N495, N499, 
        ADD_32x32_fast_I255_Y_0, N556, ADD_32x32_fast_I284_Y_0_0, 
        \un1_counter_points_snapshot[27]\, 
        ADD_32x32_fast_I263_Y_0, N580, N588, N533, 
        ADD_32x32_fast_I283_Y_0_0, 
        \un1_counter_points_snapshot[28]\, 
        ADD_32x32_fast_I126_Y_1, 
        \un1_counter_points_snapshot[20]\, N419, 
        ADD_32x32_fast_I126_Y_0, 
        \un1_counter_points_snapshot[21]\, 
        ADD_32x32_fast_I134_Y_1, 
        \un1_counter_points_snapshot[22]\, N401, 
        ADD_32x32_fast_I134_Y_0, 
        \un1_counter_points_snapshot[25]\, N404, 
        ADD_32x32_fast_I118_Y_1, N425, ADD_32x32_fast_I118_Y_0, 
        ADD_32x32_fast_I142_Y_0, 
        \un1_counter_points_snapshot_i[26]\, 
        \counter_points_snapshot_10_12_i_o2_0\, 
        un1_data_in_validlt30_28, un1_data_in_validlt30_20, 
        un1_data_in_validlt30_19, un1_data_in_validlt30_26, 
        un1_data_in_validlt30_27, un1_data_in_validlt30_16, 
        un1_data_in_validlt30_15, un1_data_in_validlt30_24, 
        un1_data_in_validlt30_12, un1_data_in_validlt30_11, 
        un1_data_in_validlt30_22, un1_data_in_validlt30_4, 
        un1_data_in_validlt30_3, un1_data_in_validlt30_18, 
        un1_data_in_validlt30_14, un1_data_in_validlt30_10, 
        \counter_points_snapshot[19]_net_1\, 
        \counter_points_snapshot[18]_net_1\, 
        un1_data_in_validlt30_8, 
        \counter_points_snapshot[14]_net_1\, 
        un1_data_in_validlt30_6, 
        \counter_points_snapshot[11]_net_1\, 
        \counter_points_snapshot[10]_net_1\, 
        un1_data_in_validlt30_2, 
        \counter_points_snapshot[3]_net_1\, 
        \counter_points_snapshot[2]_net_1\, 
        \counter_points_snapshot[1]_net_1\, 
        \counter_points_snapshot[0]_net_1\, 
        \counter_points_snapshot[28]_net_1\, 
        \counter_points_snapshot_i_0[24]\, 
        \counter_points_snapshot[23]_net_1\, 
        \counter_points_snapshot[16]_net_1\, 
        \counter_points_snapshot[17]_net_1\, 
        \counter_points_snapshot[12]_net_1\, 
        \counter_points_snapshot[8]_net_1\, 
        \counter_points_snapshot[9]_net_1\, 
        \counter_points_snapshot[6]_net_1\, 
        \counter_points_snapshot[7]_net_1\, 
        \counter_points_snapshot[4]_net_1\, 
        \counter_points_snapshot[5]_net_1\, N738, N771, N742, 
        N622, N777, \un1_data_out_valid_0_sqmuxa_2[10]\, N786, 
        \un1_data_out_valid_0_sqmuxa_2[9]\, N789_i, 
        \un1_data_out_valid_0_sqmuxa_2[5]\, N654_i, 
        \un1_data_out_valid_0_sqmuxa_2[4]\, N529, 
        \un1_data_out_valid_0_sqmuxa_2[8]\, 
        \un1_counter_points_snapshot[23]\, N648, 
        \un1_data_out_valid_0_sqmuxa_2[11]\, N783, N758, N638, 
        N740, N774, N620, N744, N752, N750, N630, N754, N634, 
        N650_i, N746, N626, N762_i, N594, N642, N764, N628, N748, 
        N766, N380, N646, N443, N440, N497, N_49, N_57, N_52, 
        N_60, counter_points_snapshot_0_sqmuxa_1, N_47, 
        \un1_data_out_valid_0_sqmuxa_2[1]\, 
        \un1_counter_points_snapshot[30]\, 
        \un1_data_out_valid_0_sqmuxa_2[2]\, 
        \un1_counter_points_snapshot_i[29]\, 
        \un1_data_out_valid_0_sqmuxa_2[6]\, N652, N756, N636, 
        N572, \un1_data_out_valid_0_sqmuxa_2[3]\, 
        \un1_data_out_valid_0_sqmuxa_2[7]\, N578, N515, N586, 
        N523, N527, N503, N570, N590, N531, N566, N582, N574, 
        N383, N768, N_20, counter_points_snapshot_2_sqmuxa_i, 
        N_21, N_25, N_26, \counter_points_snapshot_10[4]\, 
        counter_points_snapshot_2_sqmuxa_1, 
        \counter_points_snapshot_10[5]\, 
        \counter_points_snapshot_10[9]\, 
        \counter_points_snapshot_10[10]\, N_9, N_13, N_15, N_41, 
        N_45, \un1_counter_points_snapshot[31]\, 
        \counter_points_snapshot_10[0]\, N_16, 
        \un1_data_out_valid_0_sqmuxa_2[0]\, 
        \counter_points_snapshot_10[8]\, N_24, N_7, N780, 
        \counter_points_snapshot_10[11]\, N_27, N487, N_43, 
        \counter_points_snapshot_10[6]\, N_22, N422, N455, N_39, 
        N_37, N_33, N_29, \counter_points_snapshot_RNO[19]_net_1\, 
        N_35, \counter_points_snapshot_RNO[18]_net_1\, 
        \counter_points_snapshot_RNO[17]_net_1\, 
        \counter_points_snapshot_RNO[22]_net_1\, N446, N_11, N760, 
        \counter_points_snapshot_RNO[20]_net_1\, 
        \counter_points_snapshot_RNO[21]_net_1\, N_17, 
        \counter_points_snapshot_10[1]\, N386, 
        \counter_points_snapshot_10[2]\, N_18, N_31, N511, N_19, 
        \counter_points_snapshot_10[3]\, N_23, 
        \counter_points_snapshot_10[7]\, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 


    \counter_points_snapshot_RNI58FP[1]\ : MX2
      port map(A => I_5_20, B => 
        \counter_points_snapshot[1]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[30]\);
    
    \counter_points_snapshot_RNIUTOI[10]\ : NOR3A
      port map(A => un1_data_in_validlt30_6, B => 
        \counter_points_snapshot[11]_net_1\, C => 
        \counter_points_snapshot[10]_net_1\, Y => 
        un1_data_in_validlt30_18);
    
    \counter_points_snapshot[13]\ : DFN1C0
      port map(D => N_9, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[13]_net_1\);
    
    \counter_points_snapshot[11]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[11]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[11]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I284_Y_0 : AX1
      port map(A => N533, B => N529, C => 
        ADD_32x32_fast_I284_Y_0_0, Y => 
        \un1_data_out_valid_0_sqmuxa_2[4]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I26_G0N : NOR3B
      port map(A => \counter_points_snapshot[26]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N458);
    
    \data_out[110]\ : DFN1C0
      port map(D => sample_f2_wdata(46), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(110));
    
    \counter_points_snapshot_RNO_0[10]\ : MX2C
      port map(A => I_56_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[10]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_26);
    
    \counter_points_snapshot_RNO[27]\ : XA1B
      port map(A => N746, B => ADD_32x32_fast_I307_Y_0_0, C => 
        N_52, Y => N_37);
    
    \counter_points_snapshot[9]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[9]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[9]_net_1\);
    
    \counter_points_snapshot[28]\ : DFN1C0
      port map(D => N_39, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[28]_net_1\);
    
    \counter_points_snapshot_RNO[19]\ : XA1C
      port map(A => N762_i, B => ADD_32x32_fast_I299_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[19]_net_1\);
    
    \counter_points_snapshot_RNI1NC9[12]\ : NOR2
      port map(A => \counter_points_snapshot[12]_net_1\, B => 
        \counter_points_snapshot[13]_net_1\, Y => 
        un1_data_in_validlt30_6);
    
    \data_out[91]\ : DFN1C0
      port map(D => sample_f2_wdata(27), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(91));
    
    \counter_points_snapshot_RNIB9461[5]\ : MX2C
      port map(A => I_24_4, B => 
        \counter_points_snapshot[5]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot_i[26]\);
    
    \data_out[120]\ : DFN1C0
      port map(D => sample_f2_wdata(56), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(120));
    
    \counter_points_snapshot_RNO[24]\ : XO1
      port map(A => N752, B => ADD_32x32_fast_I304_Y_0_0, C => 
        N_52, Y => N_31);
    
    \counter_points_snapshot_RNIU9BB2[14]\ : NOR3C
      port map(A => un1_data_in_validlt30_20, B => 
        un1_data_in_validlt30_19, C => un1_data_in_validlt30_26, 
        Y => un1_data_in_validlt30_28);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y : NOR3
      port map(A => N626, B => ADD_32x32_fast_I254_Y_0, C => N783, 
        Y => N746);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I190_Y : OR2
      port map(A => N586, B => N578, Y => N642);
    
    \data_out[130]\ : DFN1C0
      port map(D => sample_f2_wdata(66), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(130));
    
    \data_out[104]\ : DFN1C0
      port map(D => sample_f2_wdata(40), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(104));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I104_Y : NOR3
      port map(A => N443, B => N446, C => N487, Y => N550);
    
    \counter_points_snapshot_RNO_0[4]\ : MX2C
      port map(A => I_20_12, B => 
        \un1_data_out_valid_0_sqmuxa_2[4]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_20);
    
    \counter_points_snapshot_RNO_0[1]\ : MX2C
      port map(A => I_5_20, B => 
        \un1_data_out_valid_0_sqmuxa_2[1]\, S => N_60, Y => N_17);
    
    \counter_points_snapshot_RNIJDPK[19]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[19]_net_1\, Y => 
        \un1_counter_points_snapshot[12]\);
    
    \data_out[102]\ : DFN1C0
      port map(D => sample_f2_wdata(38), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(102));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y : OR3B
      port map(A => N622, B => ADD_32x32_fast_I252_Y_1, C => N777, 
        Y => N742);
    
    \counter_points_snapshot_RNO[7]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_23, 
        Y => \counter_points_snapshot_10[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I309_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I309_Y_0_0);
    
    \counter_points_snapshot_RNO[12]\ : XA1C
      port map(A => N780, B => ADD_32x32_fast_I292_Y_0_0, C => 
        N_52, Y => N_7);
    
    \counter_points_snapshot_RNIKTDU4_0[31]\ : AO1C
      port map(A => start_snapshot_f2, B => un1_data_in_valid, C
         => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, Y => 
        N_47_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I235_Y : NOR2B
      port map(A => N650_i, B => N634, Y => N771);
    
    \data_out[93]\ : DFN1C0
      port map(D => sample_f2_wdata(29), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(93));
    
    \counter_points_snapshot[4]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[4]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[4]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I301_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[21]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I301_Y_0_0);
    
    \data_out[159]\ : DFN1C0
      port map(D => sample_f2_wdata(95), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(159));
    
    \data_out[105]\ : DFN1C0
      port map(D => sample_f2_wdata(41), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(105));
    
    \counter_points_snapshot[15]\ : DFN1C0
      port map(D => N_13, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[15]_net_1\);
    
    \data_out[141]\ : DFN1C0
      port map(D => sample_f2_wdata(77), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(141));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I108_Y : OR3
      port map(A => N443, B => N446, C => N495, Y => N554);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I140_Y : OR2A
      port map(A => N523, B => N527, Y => N586);
    
    \data_out[81]\ : DFN1C0
      port map(D => sample_f2_wdata(17), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(81));
    
    counter_points_snapshot_10_12_i_o2 : OR2B
      port map(A => \counter_points_snapshot_10_12_i_o2_0\, B => 
        N_60, Y => N_52);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I310_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I310_Y_0_0);
    
    \counter_points_snapshot[7]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[7]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[7]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y_0 : NOR3A
      port map(A => N550, B => N495, C => N499, Y => 
        ADD_32x32_fast_I256_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I234_Y_0_o2 : 
        OR2A
      port map(A => N771, B => N425, Y => N768);
    
    \data_out[114]\ : DFN1C0
      port map(D => sample_f2_wdata(50), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(114));
    
    \counter_points_snapshot[0]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[0]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[0]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I182_Y : NOR2
      port map(A => N578, B => N570, Y => N634);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I120_Y : OR3
      port map(A => N419, B => N422, C => N503, Y => N566);
    
    \counter_points_snapshot[27]\ : DFN1C0
      port map(D => N_37, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[27]_net_1\);
    
    \data_out[143]\ : DFN1C0
      port map(D => sample_f2_wdata(79), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(143));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I199_Y : NOR2B
      port map(A => N590, B => N380, Y => N654_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I110_Y : OR3
      port map(A => N443, B => N440, C => N497, Y => N556);
    
    \data_out[112]\ : DFN1C0
      port map(D => sample_f2_wdata(48), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(112));
    
    \data_out[124]\ : DFN1C0
      port map(D => sample_f2_wdata(60), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(124));
    
    \data_out[134]\ : DFN1C0
      port map(D => sample_f2_wdata(70), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(134));
    
    \counter_points_snapshot_RNIMGPV[3]\ : MX2
      port map(A => I_13_20, B => 
        \counter_points_snapshot[3]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[28]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I80_Y : AO1
      port map(A => \un1_counter_points_snapshot_i[26]\, B => 
        \un1_counter_points_snapshot[25]\, C => N_47, Y => N523);
    
    \counter_points_snapshot_RNO[28]\ : XA1B
      port map(A => N744, B => ADD_32x32_fast_I308_Y_0_0, C => 
        N_52, Y => N_39);
    
    \data_out[83]\ : DFN1C0
      port map(D => sample_f2_wdata(19), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(83));
    
    \data_out[122]\ : DFN1C0
      port map(D => sample_f2_wdata(58), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(122));
    
    \data_out[115]\ : DFN1C0
      port map(D => sample_f2_wdata(51), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(115));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I44_Y : OA1C
      port map(A => \un1_counter_points_snapshot[8]\, B => 
        \un1_counter_points_snapshot[7]\, C => N_47, Y => N487);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y_0 : AO1
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        \un1_counter_points_snapshot[17]\, C => N_47_1, Y => 
        ADD_32x32_fast_I118_Y_0);
    
    \data_out[132]\ : DFN1C0
      port map(D => sample_f2_wdata(68), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(132));
    
    \counter_points_snapshot[30]\ : DFN1C0
      port map(D => N_43, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[30]_net_1\);
    
    \data_out[96]\ : DFN1C0
      port map(D => sample_f2_wdata(32), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(96));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y : NOR3
      port map(A => N628, B => ADD_32x32_fast_I255_Y_0, C => N786, 
        Y => N748);
    
    \counter_points_snapshot_RNI20DC[2]\ : NOR3A
      port map(A => un1_data_in_validlt30_2, B => 
        \counter_points_snapshot[3]_net_1\, C => 
        \counter_points_snapshot[2]_net_1\, Y => 
        un1_data_in_validlt30_16);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I294_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[17]\, B => 
        N_47_0, Y => ADD_32x32_fast_I294_Y_0_0);
    
    \data_out[125]\ : DFN1C0
      port map(D => sample_f2_wdata(61), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(125));
    
    \data_out[135]\ : DFN1C0
      port map(D => sample_f2_wdata(71), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(135));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I15_G0N : NOR3B
      port map(A => \counter_points_snapshot[15]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N425);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0 : NOR2
      port map(A => ADD_32x32_fast_I253_Y_0_0, B => N752, Y => 
        N744);
    
    \counter_points_snapshot_RNICVG64[31]\ : AO1
      port map(A => un1_data_in_validlt30_28, B => 
        un1_data_in_validlt30_27, C => 
        \counter_points_snapshot[31]_net_1\, Y => 
        un1_data_in_valid);
    
    data_out_valid : DFN1C0
      port map(D => N_49, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        data_f2_out_valid);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I174_Y : OR3
      port map(A => N499, B => N503, C => N570, Y => N626);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I29_G0N : OR3B
      port map(A => \counter_points_snapshot[29]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        I32_un1_Y);
    
    \data_out[71]\ : DFN1C0
      port map(D => sample_f2_wdata(7), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(71));
    
    \data_out[65]\ : DFN1C0
      port map(D => sample_f2_wdata(1), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(65));
    
    \counter_points_snapshot[18]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[18]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[18]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I260_Y : OR3C
      port map(A => N638, B => N622, C => N654_i, Y => N758);
    
    \data_out[86]\ : DFN1C0
      port map(D => sample_f2_wdata(22), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(86));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I166_Y : NOR3
      port map(A => N499, B => N503, C => N554, Y => N618);
    
    \data_out[150]\ : DFN1C0
      port map(D => sample_f2_wdata(86), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(150));
    
    \counter_points_snapshot_RNINR991[6]\ : MX2C
      port map(A => I_31_5, B => 
        \counter_points_snapshot[6]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[25]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I297_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[14]\, B => 
        N_47_0, Y => ADD_32x32_fast_I297_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I296_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[15]\, B => 
        N_47_0, Y => ADD_32x32_fast_I296_Y_0_0);
    
    \data_out[148]\ : DFN1C0
      port map(D => sample_f2_wdata(84), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(148));
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I13_G0N : NOR3B
      port map(A => \counter_points_snapshot[13]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N419);
    
    \counter_points_snapshot[8]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[8]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[8]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I178_Y : OR2
      port map(A => N574, B => N566, Y => N630);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I136_Y : OR3B
      port map(A => N401, B => N523, C => N404, Y => N582);
    
    \data_out[73]\ : DFN1C0
      port map(D => sample_f2_wdata(9), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(73));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I283_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[28]\, B => 
        N_47_0, Y => ADD_32x32_fast_I283_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_3 : NOR3B
      port map(A => ADD_32x32_fast_I250_Y_1, B => N618, C => N546, 
        Y => ADD_32x32_fast_I250_Y_3);
    
    \data_out[92]\ : DFN1C0
      port map(D => sample_f2_wdata(28), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(92));
    
    \data_out[67]\ : DFN1C0
      port map(D => sample_f2_wdata(3), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(67));
    
    \data_out[107]\ : DFN1C0
      port map(D => sample_f2_wdata(43), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(107));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I14_G0N : NOR2
      port map(A => \un1_counter_points_snapshot[17]\, B => 
        N_47_1, Y => N422);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y_0 : OR3
      port map(A => N580, B => N588, C => N533, Y => 
        ADD_32x32_fast_I263_Y_0);
    
    \counter_points_snapshot_RNO[6]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_22, 
        Y => \counter_points_snapshot_10[6]\);
    
    \counter_points_snapshot_RNIQURI[26]\ : NOR3A
      port map(A => un1_data_in_validlt30_14, B => 
        \counter_points_snapshot[27]_net_1\, C => 
        \counter_points_snapshot[26]_net_1\, Y => 
        un1_data_in_validlt30_22);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I290_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[21]\, C => N786, Y => 
        \un1_data_out_valid_0_sqmuxa_2[10]\);
    
    \counter_points_snapshot[29]\ : DFN1C0
      port map(D => N_41, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[29]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I300_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I300_Y_0_0);
    
    \counter_points_snapshot_RNO[25]\ : XA1B
      port map(A => N750, B => ADD_32x32_fast_I305_Y_0_0, C => 
        N_52, Y => N_33);
    
    \counter_points_snapshot[20]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[20]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[20]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I302_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I302_Y_0_0);
    
    \counter_points_snapshot_RNIICLF1[8]\ : MX2C
      port map(A => I_45_4, B => 
        \counter_points_snapshot[8]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[23]\);
    
    \counter_points_snapshot_RNIG1PK[16]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[16]_net_1\, Y => 
        \un1_counter_points_snapshot[15]\);
    
    \counter_points_snapshot[17]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[17]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[17]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I194_Y : OR2A
      port map(A => N590, B => N582, Y => N646);
    
    \counter_points_snapshot_RNI9ND9[16]\ : NOR2
      port map(A => \counter_points_snapshot[16]_net_1\, B => 
        \counter_points_snapshot[17]_net_1\, Y => 
        un1_data_in_validlt30_8);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I88_Y : OR2A
      port map(A => N383, B => N386, Y => N531);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I292_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        N_47_0, Y => ADD_32x32_fast_I292_Y_0_0);
    
    \counter_points_snapshot_RNITFFM1[0]\ : NOR3C
      port map(A => un1_data_in_validlt30_16, B => 
        un1_data_in_validlt30_15, C => un1_data_in_validlt30_24, 
        Y => un1_data_in_validlt30_27);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y : OR2B
      port map(A => ADD_32x32_fast_I250_Y_3, B => N771, Y => N738);
    
    \data_out[154]\ : DFN1C0
      port map(D => sample_f2_wdata(90), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(154));
    
    \counter_points_snapshot_RNI047N1[11]\ : MX2
      port map(A => N_4, B => \counter_points_snapshot[11]_net_1\, 
        S => counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[20]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I261_Y_0_o2 : 
        OR2
      port map(A => N764, B => N497, Y => N760);
    
    \data_out[82]\ : DFN1C0
      port map(D => sample_f2_wdata(18), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(82));
    
    \data_out[117]\ : DFN1C0
      port map(D => sample_f2_wdata(53), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(117));
    
    \counter_points_snapshot_RNO[20]\ : XA1C
      port map(A => N760, B => ADD_32x32_fast_I300_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[20]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I254_Y_0 : OR2
      port map(A => N554, B => N546, Y => ADD_32x32_fast_I254_Y_0);
    
    \data_out[76]\ : DFN1C0
      port map(D => sample_f2_wdata(12), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(76));
    
    \data_out[152]\ : DFN1C0
      port map(D => sample_f2_wdata(88), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(152));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I118_Y_1 : OA1B
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[14]\, C => N425, Y => 
        ADD_32x32_fast_I118_Y_1);
    
    \data_out[149]\ : DFN1C0
      port map(D => sample_f2_wdata(85), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(149));
    
    \data_out[127]\ : DFN1C0
      port map(D => sample_f2_wdata(63), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(127));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I237_Y : OR2B
      port map(A => N654_i, B => N638, Y => N777);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I236_Y : NOR2
      port map(A => N652, B => N636, Y => N774);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I198_Y : OR2
      port map(A => N588, B => N533, Y => N652);
    
    \data_out[137]\ : DFN1C0
      port map(D => sample_f2_wdata(73), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(137));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I30_G0N : OR3B
      port map(A => \counter_points_snapshot[30]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N470);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I144_Y : NOR2
      port map(A => N531, B => N527, Y => N590);
    
    \data_out[155]\ : DFN1C0
      port map(D => sample_f2_wdata(91), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(155));
    
    \counter_points_snapshot_RNIV6C9[20]\ : NOR2
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        \counter_points_snapshot[21]_net_1\, Y => 
        un1_data_in_validlt30_10);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \counter_points_snapshot_RNO[5]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_21, 
        Y => \counter_points_snapshot_10[5]\);
    
    \counter_points_snapshot_RNO[17]\ : XA1C
      port map(A => N766, B => ADD_32x32_fast_I297_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[17]_net_1\);
    
    data_out_valid_RNO_0 : OR3A
      port map(A => un1_data_in_valid, B => start_snapshot_f2, C
         => burst_f2, Y => N_57);
    
    \data_out[90]\ : DFN1C0
      port map(D => sample_f2_wdata(26), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(90));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y_0 : AO1
      port map(A => \un1_counter_points_snapshot[21]\, B => 
        \un1_counter_points_snapshot[19]\, C => N_47_1, Y => 
        ADD_32x32_fast_I126_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I124_Y : OR3
      port map(A => N419, B => N422, C => N511, Y => N570);
    
    \counter_points_snapshot[2]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[2]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[2]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y : OR3B
      port map(A => ADD_32x32_fast_I251_Y_2, B => N774, C => N620, 
        Y => N740);
    
    \counter_points_snapshot_RNO[14]\ : XA1C
      port map(A => N774, B => ADD_32x32_fast_I294_Y_0_0, C => 
        N_52, Y => N_11);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I20_G0N : NOR3B
      port map(A => \counter_points_snapshot[20]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N440);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I132_Y : OR3A
      port map(A => N401, B => N404, C => N515, Y => N578);
    
    \counter_points_snapshot_RNIF7E9[28]\ : NOR2
      port map(A => \counter_points_snapshot[28]_net_1\, B => 
        \counter_points_snapshot[29]_net_1\, Y => 
        un1_data_in_validlt30_14);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I282_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot_i[29]\, C => N533, Y => 
        \un1_data_out_valid_0_sqmuxa_2[2]\);
    
    counter_points_snapshot_2_sqmuxa_0_a2 : OR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_60, 
        Y => counter_points_snapshot_2_sqmuxa_i);
    
    \data_out[99]\ : DFN1C0
      port map(D => sample_f2_wdata(35), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(99));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I258_Y : OR3C
      port map(A => N634, B => N618, C => N650_i, Y => N754);
    
    \data_out[106]\ : DFN1C0
      port map(D => sample_f2_wdata(42), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(106));
    
    \counter_points_snapshot_RNO[21]\ : XA1C
      port map(A => N758, B => ADD_32x32_fast_I301_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[21]_net_1\);
    
    \counter_points_snapshot_RNI77D9[24]\ : NOR2A
      port map(A => \counter_points_snapshot_i_0[24]\, B => 
        \counter_points_snapshot[25]_net_1\, Y => 
        un1_data_in_validlt30_12);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I128_Y : OR2
      port map(A => N515, B => N511, Y => N574);
    
    \data_out[98]\ : DFN1C0
      port map(D => sample_f2_wdata(34), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(98));
    
    \data_out[80]\ : DFN1C0
      port map(D => sample_f2_wdata(16), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(80));
    
    \data_out[72]\ : DFN1C0
      port map(D => sample_f2_wdata(8), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(72));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I256_Y : OR3B
      port map(A => ADD_32x32_fast_I256_Y_0, B => N789_i, C => 
        N630, Y => N750);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I22_G0N : NOR3B
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N446);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I56_Y : AOI1
      port map(A => \un1_counter_points_snapshot[14]\, B => 
        \un1_counter_points_snapshot[13]\, C => N_47, Y => N499);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I288_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[23]\, C => N648, Y => 
        \un1_data_out_valid_0_sqmuxa_2[8]\);
    
    counter_points_snapshot_2_sqmuxa_0_a2_0 : OR2A
      port map(A => start_snapshot_f2, B => sample_f2_val, Y => 
        N_60);
    
    \data_out[89]\ : DFN1C0
      port map(D => sample_f2_wdata(25), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(89));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I263_Y : OR2
      port map(A => ADD_32x32_fast_I263_Y_0, B => N628, Y => N764);
    
    counter_points_snapshot_0_sqmuxa_1_0_a2 : OR3B
      port map(A => sample_f2_val, B => start_snapshot_f2, C => 
        burst_f2, Y => counter_points_snapshot_0_sqmuxa_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I289_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[22]\, C => N789_i, Y => 
        \un1_data_out_valid_0_sqmuxa_2[9]\);
    
    \data_out[116]\ : DFN1C0
      port map(D => sample_f2_wdata(52), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(116));
    
    \counter_points_snapshot[19]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[19]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[19]_net_1\);
    
    \counter_points_snapshot_RNO_0[2]\ : MX2C
      port map(A => I_9_20, B => 
        \un1_data_out_valid_0_sqmuxa_2[2]\, S => N_60, Y => N_18);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I298_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[13]\, B => 
        N_47_0, Y => ADD_32x32_fast_I298_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I197_Y : NOR2
      port map(A => N594, B => N586, Y => N650_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I285_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot_i[26]\, C => N654_i, Y => 
        \un1_data_out_valid_0_sqmuxa_2[5]\);
    
    \counter_points_snapshot[10]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[10]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[10]_net_1\);
    
    \counter_points_snapshot_RNO[18]\ : XA1B
      port map(A => N764, B => ADD_32x32_fast_I298_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[18]_net_1\);
    
    \data_out[88]\ : DFN1C0
      port map(D => sample_f2_wdata(24), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(88));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_S_0 : XNOR2
      port map(A => \un1_counter_points_snapshot[31]\, B => 
        N_47_1, Y => \un1_data_out_valid_0_sqmuxa_2[0]\);
    
    \data_out[126]\ : DFN1C0
      port map(D => sample_f2_wdata(62), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(126));
    
    \data_out[94]\ : DFN1C0
      port map(D => sample_f2_wdata(30), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(94));
    
    \data_out[140]\ : DFN1C0
      port map(D => sample_f2_wdata(76), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(140));
    
    \data_out[136]\ : DFN1C0
      port map(D => sample_f2_wdata(72), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(136));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I27_G0N : OR3B
      port map(A => \counter_points_snapshot[27]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_1, Y => 
        N461);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I293_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[13]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I293_Y_0_0);
    
    \un1_data_out_valid_0_sqmuxa_1_i_0[31]\ : AOI1B
      port map(A => start_snapshot_f2, B => burst_f2, C => 
        sample_f2_val, Y => 
        \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\);
    
    \counter_points_snapshot_RNIH5PK[17]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[17]_net_1\, Y => 
        \un1_counter_points_snapshot[14]\);
    
    \counter_points_snapshot[22]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[22]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[22]_net_1\);
    
    \counter_points_snapshot_RNIEUQI[14]\ : NOR3A
      port map(A => un1_data_in_validlt30_8, B => 
        \counter_points_snapshot[15]_net_1\, C => 
        \counter_points_snapshot[14]_net_1\, Y => 
        un1_data_in_validlt30_19);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I147_Y : OR2A
      port map(A => N380, B => N531, Y => N594);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I304_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[7]\, B => N_47_0, 
        Y => ADD_32x32_fast_I304_Y_0_0);
    
    \data_out[101]\ : DFN1C0
      port map(D => sample_f2_wdata(37), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(101));
    
    \data_out[157]\ : DFN1C0
      port map(D => sample_f2_wdata(93), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(157));
    
    \counter_points_snapshot_RNO[4]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_20, 
        Y => \counter_points_snapshot_10[4]\);
    
    \counter_points_snapshot_RNO[30]\ : XA1C
      port map(A => N740, B => ADD_32x32_fast_I310_Y_0_0, C => 
        N_52, Y => N_43);
    
    \counter_points_snapshot_RNIEPOK[14]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[14]_net_1\, Y => 
        \un1_counter_points_snapshot[17]\);
    
    \counter_points_snapshot[6]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[6]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[6]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I54_Y_0_o2 : 
        AOI1
      port map(A => \un1_counter_points_snapshot[13]\, B => 
        \un1_counter_points_snapshot[12]\, C => N_47, Y => N497);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I176_Y : OR3B
      port map(A => ADD_32x32_fast_I118_Y_0, B => 
        ADD_32x32_fast_I118_Y_1, C => N572, Y => N628);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y_0 : OA1B
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[25]\, C => N404, Y => 
        ADD_32x32_fast_I134_Y_0);
    
    \data_out[70]\ : DFN1C0
      port map(D => sample_f2_wdata(6), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(70));
    
    \counter_points_snapshot_RNO_0[5]\ : MX2C
      port map(A => I_24_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[5]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_21);
    
    \data_out[84]\ : DFN1C0
      port map(D => sample_f2_wdata(20), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(84));
    
    \data_out[103]\ : DFN1C0
      port map(D => sample_f2_wdata(39), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(103));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I7_G0N : OR2A
      port map(A => \un1_counter_points_snapshot[24]\, B => N_47, 
        Y => N401);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I84_Y : OA1B
      port map(A => \un1_counter_points_snapshot[27]\, B => 
        \un1_counter_points_snapshot[28]\, C => N_47, Y => N527);
    
    \counter_points_snapshot[5]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[5]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[5]_net_1\);
    
    \counter_points_snapshot_RNO[26]\ : XA1B
      port map(A => N748, B => ADD_32x32_fast_I306_Y_0_0, C => 
        N_52, Y => N_35);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I8_G0N : NOR2
      port map(A => \un1_counter_points_snapshot[23]\, B => 
        N_47_1, Y => N404);
    
    \data_out[79]\ : DFN1C0
      port map(D => sample_f2_wdata(15), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(79));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I281_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[30]\, C => N380, Y => 
        \un1_data_out_valid_0_sqmuxa_2[1]\);
    
    \data_out[144]\ : DFN1C0
      port map(D => sample_f2_wdata(80), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(144));
    
    counter_points_snapshot_0_sqmuxa_1_0_a2_0 : OR3B
      port map(A => sample_f2_val, B => start_snapshot_f2, C => 
        burst_f2, Y => counter_points_snapshot_0_sqmuxa_1_0);
    
    \counter_points_snapshot_RNI1BRI1[9]\ : MX2C
      port map(A => I_52_4, B => 
        \counter_points_snapshot[9]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[22]\);
    
    \counter_points_snapshot_RNO[8]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_24, 
        Y => \counter_points_snapshot_10[8]\);
    
    \data_out[111]\ : DFN1C0
      port map(D => sample_f2_wdata(47), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(111));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I295_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[15]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I295_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I0_CO1 : OR2A
      port map(A => \un1_counter_points_snapshot[31]\, B => 
        N_47_1, Y => N380);
    
    \data_out[142]\ : DFN1C0
      port map(D => sample_f2_wdata(78), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(142));
    
    \data_out[78]\ : DFN1C0
      port map(D => sample_f2_wdata(14), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(78));
    
    \counter_points_snapshot_RNO[23]\ : XA1B
      port map(A => N754, B => ADD_32x32_fast_I303_Y_0_0, C => 
        N_52, Y => N_29);
    
    \counter_points_snapshot_RNIKTDU4[31]\ : AO1C
      port map(A => start_snapshot_f2, B => un1_data_in_valid, C
         => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, Y => 
        N_47_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I184_Y : OR2
      port map(A => N580, B => N572, Y => N636);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y_1 : OA1
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[22]\, C => N401, Y => 
        ADD_32x32_fast_I134_Y_1);
    
    \counter_points_snapshot_RNO_0[3]\ : MX2C
      port map(A => I_13_20, B => 
        \un1_data_out_valid_0_sqmuxa_2[3]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_19);
    
    \counter_points_snapshot[26]\ : DFN1C0
      port map(D => N_35, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[26]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I305_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[25]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I305_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I252_Y_1 : NOR3B
      port map(A => N483, B => N550, C => N479, Y => 
        ADD_32x32_fast_I252_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I1_G0N : OR2A
      port map(A => \un1_counter_points_snapshot[30]\, B => N_47, 
        Y => N383);
    
    \data_out[121]\ : DFN1C0
      port map(D => sample_f2_wdata(57), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(121));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I60_Y : AO1D
      port map(A => \un1_counter_points_snapshot[15]\, B => N_47, 
        C => N425, Y => N503);
    
    \counter_points_snapshot_RNO[0]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_16, 
        Y => \counter_points_snapshot_10[0]\);
    
    \counter_points_snapshot_RNI4IFC1[7]\ : MX2
      port map(A => I_38_4, B => 
        \counter_points_snapshot[7]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[24]\);
    
    \data_out[131]\ : DFN1C0
      port map(D => sample_f2_wdata(67), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(131));
    
    \data_out[113]\ : DFN1C0
      port map(D => sample_f2_wdata(49), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(113));
    
    \data_out[145]\ : DFN1C0
      port map(D => sample_f2_wdata(81), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(145));
    
    \data_out[66]\ : DFN1C0
      port map(D => sample_f2_wdata(2), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(66));
    
    \counter_points_snapshot[1]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[1]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[1]_net_1\);
    
    \counter_points_snapshot_RNO[31]\ : XA1B
      port map(A => N738, B => ADD_32x32_fast_I311_Y_0_0, C => 
        N_52, Y => N_45);
    
    \counter_points_snapshot_RNO_0[0]\ : MX2B
      port map(A => nb_snapshot_param(0), B => 
        \un1_data_out_valid_0_sqmuxa_2[0]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_16);
    
    \counter_points_snapshot_RNO[15]\ : XA1C
      port map(A => N771, B => ADD_32x32_fast_I295_Y_0_0, C => 
        N_52, Y => N_13);
    
    \data_out[123]\ : DFN1C0
      port map(D => sample_f2_wdata(59), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(123));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \data_out[133]\ : DFN1C0
      port map(D => sample_f2_wdata(69), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(133));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I21_G0N : NOR3B
      port map(A => \counter_points_snapshot[21]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N443);
    
    \counter_points_snapshot_RNO[29]\ : XA1C
      port map(A => N742, B => ADD_32x32_fast_I309_Y_0_0, C => 
        N_52, Y => N_41);
    
    \counter_points_snapshot[31]\ : DFN1C0
      port map(D => N_45, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[31]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I36_Y : AO1C
      port map(A => N_47_1, B => \un1_counter_points_snapshot[3]\, 
        C => N461, Y => N479);
    
    \counter_points_snapshot_RNI0RU21[4]\ : MX2
      port map(A => I_20_12, B => 
        \counter_points_snapshot[4]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[27]\);
    
    \data_out[74]\ : DFN1C0
      port map(D => sample_f2_wdata(10), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(74));
    
    \counter_points_snapshot_RNO[10]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_26, 
        Y => \counter_points_snapshot_10[10]\);
    
    \counter_points_snapshot_RNI7G66[6]\ : NOR2
      port map(A => \counter_points_snapshot[6]_net_1\, B => 
        \counter_points_snapshot[7]_net_1\, Y => 
        un1_data_in_validlt30_3);
    
    \data_out[108]\ : DFN1C0
      port map(D => sample_f2_wdata(44), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(108));
    
    \counter_points_snapshot_RNO_0[6]\ : MX2C
      port map(A => I_31_5, B => 
        \un1_data_out_valid_0_sqmuxa_2[6]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_22);
    
    \counter_points_snapshot_RNI3NC9[23]\ : NOR2
      port map(A => \counter_points_snapshot[22]_net_1\, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        un1_data_in_validlt30_11);
    
    \data_out[156]\ : DFN1C0
      port map(D => sample_f2_wdata(92), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(156));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I240_Y : OR3
      port map(A => N580, B => N588, C => N533, Y => N786);
    
    \counter_points_snapshot_RNO_0[8]\ : MX2C
      port map(A => I_45_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[8]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_24);
    
    \counter_points_snapshot_RNO[1]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_17, 
        Y => \counter_points_snapshot_10[1]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I303_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[8]\, B => N_47_0, 
        Y => ADD_32x32_fast_I303_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I25_G0N : NOR3B
      port map(A => \counter_points_snapshot[25]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1, C => N_47, Y => N455);
    
    \counter_points_snapshot_RNIGU5V[6]\ : NOR3C
      port map(A => un1_data_in_validlt30_4, B => 
        un1_data_in_validlt30_3, C => un1_data_in_validlt30_18, Y
         => un1_data_in_validlt30_24);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I40_Y : NOR2
      port map(A => N458, B => N455, Y => N483);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I257_Y_0_o2 : 
        OR2
      port map(A => N756, B => N489, Y => N752);
    
    \counter_points_snapshot_RNO[22]\ : XA1C
      port map(A => N756, B => ADD_32x32_fast_I302_Y_0_0, C => 
        N_52, Y => \counter_points_snapshot_RNO[22]_net_1\);
    
    \counter_points_snapshot[12]\ : DFN1C0
      port map(D => N_7, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[12]_net_1\);
    
    \counter_points_snapshot[24]\ : DFN1P0
      port map(D => N_31, CLK => HCLK_c, PRE => HRESETn_c, Q => 
        \counter_points_snapshot_i_0[24]\);
    
    \counter_points_snapshot_RNIKTDU4_1[31]\ : AO1C
      port map(A => start_snapshot_f2, B => un1_data_in_valid, C
         => \un1_data_out_valid_0_sqmuxa_1_i_0[31]_net_1\, Y => 
        N_47);
    
    \data_out[95]\ : DFN1C0
      port map(D => sample_f2_wdata(31), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(95));
    
    \counter_points_snapshot_RNIJ9PK[28]\ : NOR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[28]_net_1\, Y => 
        \un1_counter_points_snapshot[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I196_Y_0_o2 : 
        OR2B
      port map(A => N650_i, B => N401, Y => N648);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y : OR2B
      port map(A => ADD_32x32_fast_I126_Y_1, B => 
        ADD_32x32_fast_I126_Y_0, Y => N572);
    
    \counter_points_snapshot_RNO_0[9]\ : MX2C
      port map(A => I_52_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[9]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_25);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I126_Y_1 : OA1C
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        N_47_1, C => N419, Y => ADD_32x32_fast_I126_Y_1);
    
    \counter_points_snapshot_RNO[3]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_19, 
        Y => \counter_points_snapshot_10[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y_0 : AO1A
      port map(A => \un1_counter_points_snapshot[27]\, B => 
        \un1_counter_points_snapshot_i[26]\, C => N_47_1, Y => 
        ADD_32x32_fast_I142_Y_0);
    
    \data_out[118]\ : DFN1C0
      port map(D => sample_f2_wdata(54), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(118));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I241_Y : NOR2A
      port map(A => N380, B => N646, Y => N789_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I306_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[26]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I306_Y_0_0);
    
    \counter_points_snapshot_RNICEQI[18]\ : NOR3A
      port map(A => un1_data_in_validlt30_10, B => 
        \counter_points_snapshot[19]_net_1\, C => 
        \counter_points_snapshot[18]_net_1\, Y => 
        un1_data_in_validlt30_20);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_1 : NOR3B
      port map(A => N461, B => ADD_32x32_fast_I251_Y_0, C => N458, 
        Y => ADD_32x32_fast_I251_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I239_Y : OR2
      port map(A => N642, B => N594, Y => N783);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I287_Y_0 : XOR2
      port map(A => ADD_32x32_fast_I287_Y_0_0, B => N650_i, Y => 
        \un1_data_out_valid_0_sqmuxa_2[7]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I286_Y_0 : XOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[25]\, C => N652, Y => 
        \un1_data_out_valid_0_sqmuxa_2[6]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I46_Y_0_o2 : 
        AO1D
      port map(A => \un1_counter_points_snapshot[8]\, B => N_47, 
        C => N446, Y => N489);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I291_Y_0 : XNOR3
      port map(A => N_47_1, B => 
        \un1_counter_points_snapshot[20]\, C => N783, Y => 
        \un1_data_out_valid_0_sqmuxa_2[11]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I100_Y : OR2A
      port map(A => N483, B => N487, Y => N546);
    
    \data_out[128]\ : DFN1C0
      port map(D => sample_f2_wdata(64), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(128));
    
    \counter_points_snapshot_RNO[11]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_27, 
        Y => \counter_points_snapshot_10[11]\);
    
    \data_out[97]\ : DFN1C0
      port map(D => sample_f2_wdata(33), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(97));
    
    \data_out[138]\ : DFN1C0
      port map(D => sample_f2_wdata(74), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(138));
    
    \counter_points_snapshot_RNII9PK[18]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot[18]_net_1\, Y => 
        \un1_counter_points_snapshot[13]\);
    
    \counter_points_snapshot_RNIDAKS[2]\ : MX2C
      port map(A => I_9_20, B => 
        \counter_points_snapshot[2]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot_i[29]\);
    
    \counter_points_snapshot_RNIU9AM[0]\ : MX2A
      port map(A => nb_snapshot_param(0), B => 
        \counter_points_snapshot[0]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1_0, Y => 
        \un1_counter_points_snapshot[31]\);
    
    \data_out[85]\ : DFN1C0
      port map(D => sample_f2_wdata(21), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(85));
    
    \counter_points_snapshot[3]\ : DFN1C0
      port map(D => \counter_points_snapshot_10[3]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[3]_net_1\);
    
    \counter_points_snapshot_RNIVV6N1[10]\ : MX2C
      port map(A => I_56_4, B => 
        \counter_points_snapshot[10]_net_1\, S => 
        counter_points_snapshot_0_sqmuxa_1, Y => 
        \un1_counter_points_snapshot[21]\);
    
    \data_out[109]\ : DFN1C0
      port map(D => sample_f2_wdata(45), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(109));
    
    \counter_points_snapshot_RNI4TL51[23]\ : NOR3C
      port map(A => un1_data_in_validlt30_12, B => 
        un1_data_in_validlt30_11, C => un1_data_in_validlt30_22, 
        Y => un1_data_in_validlt30_26);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I68_Y : OA1C
      port map(A => \un1_counter_points_snapshot[19]\, B => 
        \un1_counter_points_snapshot[20]\, C => N_47, Y => N511);
    
    \counter_points_snapshot_RNIBHSA[0]\ : NOR3
      port map(A => \counter_points_snapshot[1]_net_1\, B => 
        \counter_points_snapshot[0]_net_1\, C => 
        \counter_points_snapshot[30]_net_1\, Y => 
        un1_data_in_validlt30_15);
    
    \counter_points_snapshot_RNIBG66[8]\ : NOR2
      port map(A => \counter_points_snapshot[8]_net_1\, B => 
        \counter_points_snapshot[9]_net_1\, Y => 
        un1_data_in_validlt30_4);
    
    \counter_points_snapshot[23]\ : DFN1C0
      port map(D => N_29, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[23]_net_1\);
    
    \counter_points_snapshot[21]\ : DFN1C0
      port map(D => \counter_points_snapshot_RNO[21]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[21]_net_1\);
    
    \counter_points_snapshot[16]\ : DFN1C0
      port map(D => N_15, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[16]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I255_Y_0 : OR3
      port map(A => N485, B => N489, C => N556, Y => 
        ADD_32x32_fast_I255_Y_0);
    
    \data_out[147]\ : DFN1C0
      port map(D => sample_f2_wdata(83), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(147));
    
    \data_out[151]\ : DFN1C0
      port map(D => sample_f2_wdata(87), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(151));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I299_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[12]\, B => 
        N_47_0, Y => ADD_32x32_fast_I299_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I308_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[3]\, B => N_47_0, 
        Y => ADD_32x32_fast_I308_Y_0_0);
    
    \data_out[87]\ : DFN1C0
      port map(D => sample_f2_wdata(23), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(87));
    
    counter_points_snapshot_10_12_i_o2_0 : NOR2A
      port map(A => enable_f2, B => burst_f2, Y => 
        \counter_points_snapshot_10_12_i_o2_0\);
    
    \data_out[153]\ : DFN1C0
      port map(D => sample_f2_wdata(89), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(153));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I283_Y_0 : XNOR2
      port map(A => ADD_32x32_fast_I283_Y_0_0, B => N594, Y => 
        \un1_data_out_valid_0_sqmuxa_2[3]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I259_Y : OR3
      port map(A => N636, B => N620, C => N652, Y => N756);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I86_Y : OA1C
      port map(A => \un1_counter_points_snapshot[28]\, B => N_47, 
        C => N386, Y => N529);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I142_Y : OR2B
      port map(A => ADD_32x32_fast_I142_Y_0, B => N529, Y => N588);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I307_Y_0_0 : 
        AX1C
      port map(A => \counter_points_snapshot[27]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I307_Y_0_0);
    
    \data_out[119]\ : DFN1C0
      port map(D => sample_f2_wdata(55), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(119));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I250_Y_1 : NOR3B
      port map(A => I32_un1_Y, B => N470, C => N479, Y => 
        ADD_32x32_fast_I250_Y_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I72_Y : AOI1
      port map(A => \un1_counter_points_snapshot[22]\, B => 
        \un1_counter_points_snapshot[21]\, C => N_47, Y => N515);
    
    \counter_points_snapshot_RNIELOK[23]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1_0, B => 
        \counter_points_snapshot[23]_net_1\, Y => 
        \un1_counter_points_snapshot[8]\);
    
    \counter_points_snapshot_RNO_0[7]\ : MX2C
      port map(A => I_38_4, B => 
        \un1_data_out_valid_0_sqmuxa_2[7]\, S => 
        counter_points_snapshot_2_sqmuxa_i, Y => N_23);
    
    \counter_points_snapshot_RNO[9]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_25, 
        Y => \counter_points_snapshot_10[9]\);
    
    \counter_points_snapshot_RNIFPOK[24]\ : NOR2A
      port map(A => counter_points_snapshot_0_sqmuxa_1, B => 
        \counter_points_snapshot_i_0[24]\, Y => 
        \un1_counter_points_snapshot[7]\);
    
    \data_out[69]\ : DFN1C0
      port map(D => sample_f2_wdata(5), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(69));
    
    \data_out[129]\ : DFN1C0
      port map(D => sample_f2_wdata(65), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(129));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I311_Y_0_0 : 
        AX1E
      port map(A => \counter_points_snapshot[31]_net_1\, B => 
        counter_points_snapshot_0_sqmuxa_1_0, C => N_47_0, Y => 
        ADD_32x32_fast_I311_Y_0_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_2 : NOR3A
      port map(A => ADD_32x32_fast_I251_Y_1, B => N485, C => N489, 
        Y => ADD_32x32_fast_I251_Y_2);
    
    \data_out[139]\ : DFN1C0
      port map(D => sample_f2_wdata(75), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(139));
    
    \counter_points_snapshot[25]\ : DFN1C0
      port map(D => N_33, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[25]_net_1\);
    
    counter_points_snapshot_2_sqmuxa_0_a2_1 : OR2A
      port map(A => enable_f2, B => burst_f2, Y => 
        counter_points_snapshot_2_sqmuxa_1);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I134_Y : OR2B
      port map(A => ADD_32x32_fast_I134_Y_1, B => 
        ADD_32x32_fast_I134_Y_0, Y => N580);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I238_Y_0_o2 : 
        OA1C
      port map(A => \un1_counter_points_snapshot[20]\, B => 
        N_47_1, C => N783, Y => N780);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I90_Y : OR2B
      port map(A => N383, B => N380, Y => N533);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I42_Y : AO1A
      port map(A => N_47, B => \un1_counter_points_snapshot[7]\, 
        C => N455, Y => N485);
    
    \data_out[75]\ : DFN1C0
      port map(D => sample_f2_wdata(11), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(75));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I284_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[27]\, B => 
        N_47_0, Y => ADD_32x32_fast_I284_Y_0_0);
    
    \data_out[68]\ : DFN1C0
      port map(D => sample_f2_wdata(4), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(68));
    
    \counter_points_snapshot_RNICHOK[12]\ : OR2B
      port map(A => counter_points_snapshot_0_sqmuxa_1_0, B => 
        \counter_points_snapshot[12]_net_1\, Y => 
        \un1_counter_points_snapshot[19]\);
    
    \counter_points_snapshot_RNI3G66[4]\ : NOR2
      port map(A => \counter_points_snapshot[4]_net_1\, B => 
        \counter_points_snapshot[5]_net_1\, Y => 
        un1_data_in_validlt30_2);
    
    \counter_points_snapshot_RNO_0[11]\ : MX2C
      port map(A => N_4, B => \un1_data_out_valid_0_sqmuxa_2[11]\, 
        S => counter_points_snapshot_2_sqmuxa_i, Y => N_27);
    
    \counter_points_snapshot[14]\ : DFN1C0
      port map(D => N_11, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \counter_points_snapshot[14]_net_1\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I251_Y_0 : OA1A
      port map(A => \un1_counter_points_snapshot[3]\, B => N_47_0, 
        C => I32_un1_Y, Y => ADD_32x32_fast_I251_Y_0);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I52_Y : AO1D
      port map(A => \un1_counter_points_snapshot[12]\, B => N_47, 
        C => N440, Y => N495);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I168_Y : OR3B
      port map(A => ADD_32x32_fast_I118_Y_0, B => 
        ADD_32x32_fast_I118_Y_1, C => N556, Y => N620);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I264_Y : NOR3A
      port map(A => N380, B => N646, C => N630, Y => N766);
    
    \counter_points_snapshot_RNO[16]\ : XA1B
      port map(A => N768, B => ADD_32x32_fast_I296_Y_0_0, C => 
        N_52, Y => N_15);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I170_Y : NOR3
      port map(A => N495, B => N499, C => N566, Y => N622);
    
    data_out_valid_RNO : NOR3C
      port map(A => sample_f2_val, B => enable_f2, C => N_57, Y
         => N_49);
    
    \data_out[100]\ : DFN1C0
      port map(D => sample_f2_wdata(36), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(100));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I262_Y : NOR3
      port map(A => N626, B => N594, C => N642, Y => N762_i);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I253_Y_0_0 : 
        OR3A
      port map(A => N461, B => N458, C => N485, Y => 
        ADD_32x32_fast_I253_Y_0_0);
    
    \data_out[77]\ : DFN1C0
      port map(D => sample_f2_wdata(13), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(77));
    
    \data_out[146]\ : DFN1C0
      port map(D => sample_f2_wdata(82), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(146));
    
    \counter_points_snapshot_RNO[2]\ : NOR2
      port map(A => counter_points_snapshot_2_sqmuxa_1, B => N_18, 
        Y => \counter_points_snapshot_10[2]\);
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I186_Y : NOR2
      port map(A => N582, B => N574, Y => N638);
    
    \counter_points_snapshot_RNO[13]\ : XA1B
      port map(A => N777, B => ADD_32x32_fast_I293_Y_0_0, C => 
        N_52, Y => N_9);
    
    \data_out[158]\ : DFN1C0
      port map(D => sample_f2_wdata(94), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(158));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I2_G0N : NOR2
      port map(A => \un1_counter_points_snapshot_i[29]\, B => 
        N_47, Y => N386);
    
    \data_out[64]\ : DFN1C0
      port map(D => sample_f2_wdata(0), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => data_f2_out(64));
    
    un1_data_out_valid_0_sqmuxa_2_ADD_32x32_fast_I287_Y_0_0 : 
        XOR2
      port map(A => \un1_counter_points_snapshot[24]\, B => 
        N_47_0, Y => ADD_32x32_fast_I287_Y_0_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\ is

    port( nb_burst_available  : in    std_logic_vector(10 downto 0);
          status_full_err     : out   std_logic_vector(2 to 2);
          status_full         : out   std_logic_vector(2 to 2);
          sel_data            : in    std_logic_vector(1 to 1);
          sel_data_1          : in    std_logic_vector(1 to 1);
          sel_data_0          : in    std_logic_vector(1 to 1);
          update_and_sel_3    : in    std_logic_vector(5 downto 4);
          addr_data_f2        : in    std_logic_vector(31 downto 0);
          status_full_ack     : in    std_logic_vector(2 to 2);
          addr_data_vector_62 : out   std_logic;
          addr_data_vector_61 : out   std_logic;
          addr_data_vector_5  : in    std_logic;
          addr_data_vector_4  : in    std_logic;
          addr_data_vector_3  : in    std_logic;
          addr_data_vector_0  : in    std_logic;
          addr_data_vector_12 : in    std_logic;
          addr_data_vector_11 : in    std_logic;
          addr_data_vector_9  : in    std_logic;
          addr_data_vector_7  : in    std_logic;
          addr_data_vector_6  : in    std_logic;
          addr_data_vector_26 : in    std_logic;
          addr_data_vector_24 : in    std_logic;
          addr_data_vector_22 : in    std_logic;
          addr_data_vector_28 : in    std_logic;
          addr_data_vector_66 : out   std_logic;
          addr_data_vector_65 : out   std_logic;
          addr_data_vector_91 : out   std_logic;
          addr_data_vector_89 : out   std_logic;
          addr_data_vector_87 : out   std_logic;
          addr_data_vector_63 : out   std_logic;
          addr_data_vector_72 : out   std_logic;
          addr_data_vector_74 : out   std_logic;
          addr_data_vector_79 : out   std_logic;
          addr_data_vector_78 : out   std_logic;
          addr_data_vector_81 : out   std_logic;
          addr_data_vector_80 : out   std_logic;
          addr_data_vector_84 : out   std_logic;
          addr_data_vector_85 : out   std_logic;
          addr_data_vector_77 : out   std_logic;
          addr_data_vector_82 : out   std_logic;
          addr_data_vector_83 : out   std_logic;
          N_1329              : out   std_logic;
          N_1328              : out   std_logic;
          N_1327              : out   std_logic;
          N_1324              : out   std_logic;
          N_1322              : out   std_logic;
          N_1321              : out   std_logic;
          N_1319              : out   std_logic;
          N_1317              : out   std_logic;
          N_1316              : out   std_logic;
          N_1308              : out   std_logic;
          N_1306              : out   std_logic;
          N_1304              : out   std_logic;
          N_1296              : out   std_logic;
          HRESETn_c           : in    std_logic;
          HCLK_c              : in    std_logic
        );

end 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\ is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \state_0[0]_net_1\, N_118, N_38, \nb_send[1]_net_1\, 
        \nb_send[0]_net_1\, N_30, \nb_send[3]_net_1\, 
        \DWACT_FINC_E[0]\, N_7, \nb_send[8]_net_1\, 
        \DWACT_FINC_E[4]\, m41_m6_0_a2_7, m41_m6_0_a2_2, 
        m41_m6_0_a2_1, m41_m6_0_a2_6, m41_m6_0_a2_4, 
        m26_m6_0_a2_6, \addr_data_vector[76]\, m26_m6_0_a2_4, 
        m26_m6_0_a2_5, \addr_data_vector[73]\, 
        \addr_data_vector[72]\, m26_m6_0_a2_2, 
        \addr_data_vector[71]\, \addr_data_vector[79]\, 
        \addr_data_vector[78]\, \addr_data_vector[74]\, 
        \un1_state_12_3_0[4]\, \update_r_i[0]\, 
        \update_r[1]_net_1\, \state_ns_i_0[3]\, N_131, 
        \un1_state_12[4]\, \un1_state_12_2[4]\, \un1_address[6]\, 
        address_0_sqmuxa, \addr_data_vector[70]\, N_5_0, N_116, 
        N_129, \state[1]_net_1\, \state_ns[0]\, N_125, N_124, 
        N_110, \state[3]_net_1\, \state[4]_net_1\, N_130, 
        \state[2]_net_1\, state7, un3_update_r, N_27_0_i_0, 
        N_13_0, N_15_0_i_0, N_16_0, N_17_0_i_0, N_19_0, 
        N_20_0_i_0, \addr_data_vector[75]\, N_22_0_i_0, N_23_0, 
        N_26_0_i_0, N_25_0, N_28_0_i_0, \addr_data_vector[80]\, 
        N_30_0_i_0, \addr_data_vector[81]\, N_31_0, 
        \un1_address[19]\, \addr_data_vector[82]\, 
        \addr_data_vector[83]\, N_34_0, \un1_address[20]\, 
        \addr_data_vector[84]\, N_37_0, \addr_data_vector[85]\, 
        \un1_address[23]\, \addr_data_vector[86]\, 
        \addr_data_vector[87]\, N_40_i_0, N_41, N_43, 
        \addr_data_vector[89]\, N_45, \addr_data_vector[91]\, 
        N_47, \addr_data_vector[93]\, N_49_i_0, 
        \addr_data_vector[95]\, N_50_i_0, \addr_data_vector[66]\, 
        \addr_data_vector[67]\, N_51_i_0, N_69, N_52_i_0, 
        \addr_data_vector[68]\, N_1_i_0, N_54_0_i_0, N_55_0_i_0, 
        \addr_data_vector[77]\, \un1_address[18]\, 
        \un1_address[21]\, \un1_address[22]\, \un1_address[24]\, 
        \addr_data_vector[88]\, \un1_address[25]\, 
        \un1_address[26]\, \addr_data_vector[90]\, 
        \un1_address[27]\, \un1_address[28]\, 
        \addr_data_vector[92]\, \un1_address[29]\, 
        \un1_address[30]\, \addr_data_vector[94]\, 
        \addr_data_vector[69]\, \address_7[2]\, \address_7[3]\, 
        \address_7[4]\, \address_7[5]\, \address_7[6]\, 
        \address_7[7]\, \address_7[8]\, \address_7[9]\, 
        \address_7[10]\, \address_7[11]\, \address_7[12]\, 
        \address_7[13]\, \address_7[15]\, \address_7[16]\, 
        \address_7[17]\, \address_7[18]\, \address_7[19]\, 
        \state[0]_net_1\, \address_7[20]\, \address_7[21]\, 
        \address_7[22]\, \address_7[23]\, \address_7[24]\, 
        \address_7[25]\, \address_7[26]\, \address_7[27]\, 
        \address_7[28]\, \address_7[29]\, \address_7[30]\, 
        \address_7[31]\, N_56_0_i_0, un1_state_9, \nb_send_5[0]\, 
        \nb_send_5[1]\, \un2_nb_send_next[1]\, \nb_send_5[2]\, 
        \un2_nb_send_next[2]\, \nb_send_5[3]\, 
        \un2_nb_send_next[3]\, \nb_send_5[4]\, 
        \un2_nb_send_next[4]\, \nb_send_5[5]\, 
        \un2_nb_send_next[5]\, \nb_send_5[6]\, 
        \un2_nb_send_next[6]\, \nb_send_5[7]\, 
        \un2_nb_send_next[7]\, \nb_send_5[8]\, 
        \un2_nb_send_next[8]\, \nb_send_5[9]\, 
        \un2_nb_send_next[9]\, \nb_send_5[10]\, 
        \un2_nb_send_next[10]\, N_126, N_113, \state_ns[2]\, 
        un1_state_11, \address_7[14]\, \nb_send[2]_net_1\, 
        \nb_send[4]_net_1\, \nb_send[5]_net_1\, 
        \nb_send[6]_net_1\, \nb_send[7]_net_1\, 
        \nb_send[9]_net_1\, \nb_send[10]_net_1\, N_4, 
        \DWACT_FINC_E[2]\, \DWACT_FINC_E[3]\, N_12, N_17, N_22, 
        \DWACT_FINC_E[1]\, N_27, N_35, \DWACT_COMP0_E[1]\, 
        \DWACT_COMP0_E[2]\, \DWACT_COMP0_E[0]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, \ACT_LT4_E[3]\, 
        \ACT_LT4_E[6]\, \ACT_LT4_E[10]\, \ACT_LT4_E[7]\, 
        \ACT_LT4_E[8]\, \ACT_LT4_E[5]\, \ACT_LT4_E[4]\, 
        \ACT_LT4_E[0]\, \ACT_LT4_E[1]\, \ACT_LT4_E[2]\, 
        \ACT_LT2_E[0]\, \ACT_LT2_E[1]\, \ACT_LT2_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, N_37, 
        N_36, N_35_0, N_32, N_34, N_33, N_31, N_28, N_29, N_30_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, 
        \DWACT_BL_EQUAL_0_E[4]\, \DWACT_BL_EQUAL_0_E[3]\, 
        \DWACT_BL_EQUAL_0_E_0[0]\, \DWACT_BL_EQUAL_0_E_0[1]\, 
        \DWACT_BL_EQUAL_0_E[2]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    addr_data_vector_66 <= \addr_data_vector[69]\;
    addr_data_vector_65 <= \addr_data_vector[68]\;
    addr_data_vector_91 <= \addr_data_vector[94]\;
    addr_data_vector_89 <= \addr_data_vector[92]\;
    addr_data_vector_87 <= \addr_data_vector[90]\;
    addr_data_vector_63 <= \addr_data_vector[66]\;
    addr_data_vector_72 <= \addr_data_vector[75]\;
    addr_data_vector_74 <= \addr_data_vector[77]\;
    addr_data_vector_79 <= \addr_data_vector[82]\;
    addr_data_vector_78 <= \addr_data_vector[81]\;
    addr_data_vector_81 <= \addr_data_vector[84]\;
    addr_data_vector_80 <= \addr_data_vector[83]\;
    addr_data_vector_84 <= \addr_data_vector[87]\;
    addr_data_vector_85 <= \addr_data_vector[88]\;
    addr_data_vector_77 <= \addr_data_vector[80]\;
    addr_data_vector_82 <= \addr_data_vector[85]\;
    addr_data_vector_83 <= \addr_data_vector[86]\;

    \address[16]\ : DFN1C0
      port map(D => \address_7[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[80]\);
    
    \address[10]\ : DFN1C0
      port map(D => \address_7[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[74]\);
    
    \state[0]\ : DFN1C0
      port map(D => N_118, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[0]_net_1\);
    
    \address[30]\ : DFN1C0
      port map(D => \address_7[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[94]\);
    
    \address_RNO[26]\ : MX2
      port map(A => \un1_address[26]\, B => addr_data_f2(26), S
         => \state[0]_net_1\, Y => \address_7[26]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_25\ : AO1C
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_31, Y => N_36);
    
    un1_address_m61 : XOR2
      port map(A => N_43, B => \addr_data_vector[90]\, Y => 
        \un1_address[26]\);
    
    \address_RNILG94[25]\ : MX2C
      port map(A => addr_data_vector_22, B => 
        \addr_data_vector[89]\, S => sel_data_1(1), Y => N_1304);
    
    \address[26]\ : DFN1C0
      port map(D => \address_7[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[90]\);
    
    \address[20]\ : DFN1C0
      port map(D => \address_7[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[84]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_42\ : AO1C
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => \un2_nb_send_next[5]\, Y => 
        \ACT_LT2_E[1]\);
    
    \address_RNI5894[10]\ : MX2C
      port map(A => addr_data_vector_7, B => 
        \addr_data_vector[74]\, S => sel_data_1(1), Y => N_1317);
    
    \FSM_SELECT_ADDRESS.state7_0_I_57\ : NOR2A
      port map(A => \ACT_LT4_E[4]\, B => \ACT_LT4_E[5]\, Y => 
        \ACT_LT4_E[6]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_36\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[1]\, B => 
        \DWACT_BL_EQUAL_0_E[0]\, Y => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\);
    
    un1_address_m51 : AX1C
      port map(A => \addr_data_vector[68]\, B => N_69, C => 
        \addr_data_vector[69]\, Y => N_52_i_0);
    
    un1_address_m26_m6_0_a2_6 : NOR3C
      port map(A => \addr_data_vector[77]\, B => 
        \addr_data_vector[76]\, C => m26_m6_0_a2_4, Y => 
        m26_m6_0_a2_6);
    
    \address[12]\ : DFN1C0
      port map(D => \address_7[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[76]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_22\ : OA1A
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_29, Y => N_33);
    
    un1_address_m26_m6_0_a2 : OR3B
      port map(A => m26_m6_0_a2_6, B => m26_m6_0_a2_5, C => 
        N_13_0, Y => N_27_0_i_0);
    
    \address_RNO[29]\ : MX2
      port map(A => \un1_address[29]\, B => addr_data_f2(29), S
         => \state[0]_net_1\, Y => \address_7[29]\);
    
    un1_address_m41_m6_0_a2_7 : NOR3C
      port map(A => m41_m6_0_a2_2, B => m41_m6_0_a2_1, C => 
        m41_m6_0_a2_6, Y => m41_m6_0_a2_7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_8\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, B => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, Y => 
        \DWACT_COMP0_E[1]\);
    
    un1_address_m19 : XNOR2
      port map(A => N_19_0, B => \addr_data_vector[75]\, Y => 
        N_20_0_i_0);
    
    \address[22]\ : DFN1C0
      port map(D => \address_7[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[86]\);
    
    \address_RNO[23]\ : MX2
      port map(A => \un1_address[23]\, B => addr_data_f2(23), S
         => \state[0]_net_1\, Y => \address_7[23]\);
    
    \address[2]\ : DFN1C0
      port map(D => \address_7[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[66]\);
    
    un2_nb_send_next_I_13 : XOR2
      port map(A => N_35, B => \nb_send[3]_net_1\, Y => 
        \un2_nb_send_next[3]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_54\ : AOI1A
      port map(A => \ACT_LT4_E[0]\, B => \ACT_LT4_E[1]\, C => 
        \ACT_LT4_E[2]\, Y => \ACT_LT4_E[3]\);
    
    \address_RNO[24]\ : MX2
      port map(A => \un1_address[24]\, B => addr_data_f2(24), S
         => \state[0]_net_1\, Y => \address_7[24]\);
    
    \address_RNO[10]\ : MX2
      port map(A => N_54_0_i_0, B => addr_data_f2(10), S => 
        \state_0[0]_net_1\, Y => \address_7[10]\);
    
    \status_full_err\ : DFN1E0C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_110, Q => status_full_err(2));
    
    un2_nb_send_next_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \nb_send[8]_net_1\, C
         => \nb_send[9]_net_1\, Y => N_4);
    
    un1_address_m18 : OR3B
      port map(A => \addr_data_vector[73]\, B => 
        \addr_data_vector[74]\, C => N_16_0, Y => N_19_0);
    
    \nb_send_RNO[1]\ : NOR2B
      port map(A => \un2_nb_send_next[1]\, B => state7, Y => 
        \nb_send_5[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_51\ : NOR2B
      port map(A => \nb_send[0]_net_1\, B => 
        nb_burst_available(0), Y => \ACT_LT4_E[0]\);
    
    \address_RNIPNMA[3]\ : MX2C
      port map(A => addr_data_vector_0, B => 
        \addr_data_vector[67]\, S => sel_data_1(1), Y => N_1324);
    
    un2_nb_send_next_I_31 : XOR2
      port map(A => N_22, B => \nb_send[6]_net_1\, Y => 
        \un2_nb_send_next[6]\);
    
    \nb_send[9]\ : DFN1E0C0
      port map(D => \nb_send_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[9]_net_1\);
    
    \address_RNO[9]\ : MX2
      port map(A => N_17_0_i_0, B => addr_data_f2(9), S => 
        \state_0[0]_net_1\, Y => \address_7[9]\);
    
    \address[5]\ : DFN1C0
      port map(D => \address_7[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[69]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_5\ : XNOR2
      port map(A => \un2_nb_send_next[7]\, B => 
        nb_burst_available(7), Y => \DWACT_BL_EQUAL_0_E_0[1]\);
    
    \address[15]\ : DFN1C0
      port map(D => \address_7[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[79]\);
    
    \address[13]\ : DFN1C0
      port map(D => \address_7[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[77]\);
    
    \state[4]\ : DFN1P0
      port map(D => \state_ns[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[4]_net_1\);
    
    \nb_send_RNO[9]\ : NOR2B
      port map(A => \un2_nb_send_next[9]\, B => state7, Y => 
        \nb_send_5[9]\);
    
    \address[19]\ : DFN1C0
      port map(D => \address_7[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[83]\);
    
    \address[25]\ : DFN1C0
      port map(D => \address_7[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[89]\);
    
    \address_RNIT9IB[7]\ : MX2C
      port map(A => addr_data_vector_4, B => 
        \addr_data_vector[71]\, S => sel_data(1), Y => N_1328);
    
    un2_nb_send_next_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => \nb_send[5]_net_1\, Y => N_22);
    
    \state_RNIV5SU8[3]\ : OR3B
      port map(A => \state[3]_net_1\, B => state7, C => 
        un3_update_r, Y => address_0_sqmuxa);
    
    \address_RNIR1IB[6]\ : MX2C
      port map(A => addr_data_vector_3, B => 
        \addr_data_vector[70]\, S => sel_data(1), Y => N_1327);
    
    \address[23]\ : DFN1C0
      port map(D => \address_7[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[87]\);
    
    un1_address_m26_m6_0_a2_5 : NOR3C
      port map(A => \addr_data_vector[73]\, B => 
        \addr_data_vector[72]\, C => m26_m6_0_a2_2, Y => 
        m26_m6_0_a2_5);
    
    \state_RNISHSP8_0[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => state7, Y => N_126);
    
    un1_address_m14 : AX1
      port map(A => N_13_0, B => \addr_data_vector[71]\, C => 
        \addr_data_vector[72]\, Y => N_15_0_i_0);
    
    un1_address_m29 : AX1
      port map(A => N_27_0_i_0, B => \addr_data_vector[80]\, C
         => \addr_data_vector[81]\, Y => N_30_0_i_0);
    
    un2_nb_send_next_I_12 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => N_35);
    
    \FSM_SELECT_ADDRESS.state7_0_I_19\ : NOR2A
      port map(A => nb_burst_available(6), B => 
        \un2_nb_send_next[6]\, Y => N_30_0);
    
    \address[29]\ : DFN1C0
      port map(D => \address_7[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[93]\);
    
    \address[18]\ : DFN1C0
      port map(D => \address_7[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[82]\);
    
    \nb_send_RNO[6]\ : NOR2B
      port map(A => \un2_nb_send_next[6]\, B => state7, Y => 
        \nb_send_5[6]\);
    
    \address_RNO[21]\ : MX2
      port map(A => \un1_address[21]\, B => addr_data_f2(21), S
         => \state[0]_net_1\, Y => \address_7[21]\);
    
    \address_RNO[16]\ : MX2
      port map(A => N_28_0_i_0, B => addr_data_f2(16), S => 
        \state_0[0]_net_1\, Y => \address_7[16]\);
    
    un2_nb_send_next_I_51 : NOR2B
      port map(A => \nb_send[8]_net_1\, B => \DWACT_FINC_E[4]\, Y
         => N_7);
    
    \address[0]\ : DFN1E1C0
      port map(D => addr_data_f2(0), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        addr_data_vector_61);
    
    \address_RNITG94[29]\ : MX2C
      port map(A => addr_data_vector_26, B => 
        \addr_data_vector[93]\, S => sel_data_1(1), Y => N_1308);
    
    \state_RNIV5SU8_0[3]\ : AO1B
      port map(A => un3_update_r, B => state7, C => 
        \state[3]_net_1\, Y => un1_state_9);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \address_RNO[27]\ : MX2
      port map(A => \un1_address[27]\, B => addr_data_f2(27), S
         => \state[0]_net_1\, Y => \address_7[27]\);
    
    \address[4]\ : DFN1C0
      port map(D => \address_7[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[68]\);
    
    \address[28]\ : DFN1C0
      port map(D => \address_7[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[92]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_7\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[4]\, B => 
        \DWACT_BL_EQUAL_0_E[3]\, Y => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\);
    
    \nb_send_RNO[2]\ : NOR2B
      port map(A => \un2_nb_send_next[2]\, B => state7, Y => 
        \nb_send_5[2]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \state_RNO_0[4]\ : OR3B
      port map(A => N_131, B => N_129, C => \state[3]_net_1\, Y
         => N_125);
    
    \address_RNI9894[12]\ : MX2C
      port map(A => addr_data_vector_9, B => 
        \addr_data_vector[76]\, S => sel_data_1(1), Y => N_1319);
    
    \FSM_SELECT_ADDRESS.state7_0_I_58\ : NOR2A
      port map(A => \un2_nb_send_next[2]\, B => 
        nb_burst_available(2), Y => \ACT_LT4_E[7]\);
    
    \nb_send_RNO[7]\ : NOR2B
      port map(A => \un2_nb_send_next[7]\, B => state7, Y => 
        \nb_send_5[7]\);
    
    un2_nb_send_next_I_24 : XOR2
      port map(A => N_27, B => \nb_send[5]_net_1\, Y => 
        \un2_nb_send_next[5]\);
    
    un2_nb_send_next_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \nb_send[3]_net_1\, C
         => \nb_send[4]_net_1\, Y => N_27);
    
    un1_address_ADD_32x32_fast_I164_Y_0 : XOR3
      port map(A => address_0_sqmuxa, B => \addr_data_vector[70]\, 
        C => N_5_0, Y => \un1_address[6]\);
    
    \address_RNO[19]\ : MX2
      port map(A => \un1_address[19]\, B => addr_data_f2(19), S
         => \state[0]_net_1\, Y => \address_7[19]\);
    
    un1_address_m24 : OR3B
      port map(A => \addr_data_vector[77]\, B => 
        \addr_data_vector[78]\, C => N_23_0, Y => N_25_0);
    
    \nb_send[7]\ : DFN1E0C0
      port map(D => \nb_send_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[7]_net_1\);
    
    \update_r_RNIV5SU8[0]\ : NOR2
      port map(A => \un1_state_12_3_0[4]\, B => 
        \un1_state_12_2[4]\, Y => \un1_state_12[4]\);
    
    \address_RNO[13]\ : MX2
      port map(A => N_55_0_i_0, B => addr_data_f2(13), S => 
        \state_0[0]_net_1\, Y => \address_7[13]\);
    
    \address[14]\ : DFN1C0
      port map(D => \address_7[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[78]\);
    
    \state_RNO[1]\ : OA1C
      port map(A => N_129, B => \state[1]_net_1\, C => 
        \state_ns_i_0[3]\, Y => N_116);
    
    \nb_send[0]\ : DFN1E0C0
      port map(D => \nb_send_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[0]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_53\ : AND2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[2]\);
    
    \nb_send[6]\ : DFN1E0C0
      port map(D => \nb_send_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[6]_net_1\);
    
    \nb_send[10]\ : DFN1E0C0
      port map(D => \nb_send_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[10]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_56\ : NOR2A
      port map(A => nb_burst_available(3), B => 
        \un2_nb_send_next[3]\, Y => \ACT_LT4_E[5]\);
    
    \address_RNO[14]\ : MX2
      port map(A => N_56_0_i_0, B => addr_data_f2(14), S => 
        \state[0]_net_1\, Y => \address_7[14]\);
    
    \address_RNIPG94[27]\ : MX2C
      port map(A => addr_data_vector_24, B => 
        \addr_data_vector[91]\, S => sel_data_1(1), Y => N_1306);
    
    \nb_send_RNO[3]\ : NOR2B
      port map(A => \un2_nb_send_next[3]\, B => state7, Y => 
        \nb_send_5[3]\);
    
    \nb_send[2]\ : DFN1E0C0
      port map(D => \nb_send_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[2]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_27\ : OA1
      port map(A => N_37, B => N_36, C => N_35_0, Y => 
        \DWACT_COMP0_E[0]\);
    
    \address[24]\ : DFN1C0
      port map(D => \address_7[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[88]\);
    
    un1_address_m27 : XNOR2
      port map(A => N_27_0_i_0, B => \addr_data_vector[80]\, Y
         => N_28_0_i_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un1_address_m60 : AX1
      port map(A => N_27_0_i_0, B => m41_m6_0_a2_7, C => 
        \addr_data_vector[89]\, Y => \un1_address[25]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_44\ : AND3A
      port map(A => \ACT_LT2_E[0]\, B => \ACT_LT2_E[1]\, C => 
        \ACT_LT2_E[2]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\);
    
    un1_address_m30 : OR3B
      port map(A => \addr_data_vector[80]\, B => 
        \addr_data_vector[81]\, C => N_27_0_i_0, Y => N_31_0);
    
    \nb_send[4]\ : DFN1E0C0
      port map(D => \nb_send_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[4]_net_1\);
    
    un1_address_m16 : XNOR2
      port map(A => N_16_0, B => \addr_data_vector[73]\, Y => 
        N_17_0_i_0);
    
    un2_nb_send_next_I_45 : XOR2
      port map(A => N_12, B => \nb_send[8]_net_1\, Y => 
        \un2_nb_send_next[8]\);
    
    \nb_send_RNO[0]\ : NOR2A
      port map(A => state7, B => \nb_send[0]_net_1\, Y => 
        \nb_send_5[0]\);
    
    \nb_send_RNO[8]\ : NOR2B
      port map(A => \un2_nb_send_next[8]\, B => state7, Y => 
        \nb_send_5[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_41\ : AND2A
      port map(A => nb_burst_available(5), B => 
        \un2_nb_send_next[5]\, Y => \ACT_LT2_E[0]\);
    
    \state_RNO[4]\ : OR3C
      port map(A => N_125, B => N_124, C => \un1_state_12_2[4]\, 
        Y => \state_ns[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_4\ : XNOR2
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), Y => \DWACT_BL_EQUAL_0_E[3]\);
    
    \address[8]\ : DFN1C0
      port map(D => \address_7[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[72]\);
    
    un1_address_m50 : XOR2
      port map(A => N_69, B => \addr_data_vector[68]\, Y => 
        N_51_i_0);
    
    un1_address_m39 : XOR2
      port map(A => \un1_state_12[4]\, B => 
        \addr_data_vector[66]\, Y => N_40_i_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_24\ : OR2A
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => N_35_0);
    
    \state_ns_i_a2[1]\ : NOR2A
      port map(A => update_and_sel_3(4), B => update_and_sel_3(5), 
        Y => N_129);
    
    \address_RNO[6]\ : MX2
      port map(A => \un1_address[6]\, B => addr_data_f2(6), S => 
        \state_0[0]_net_1\, Y => \address_7[6]\);
    
    \state_RNO[2]\ : AO1A
      port map(A => status_full_ack(2), B => N_130, C => N_126, Y
         => \state_ns[2]\);
    
    \address_RNO[28]\ : MX2
      port map(A => \un1_address[28]\, B => addr_data_f2(28), S
         => \state[0]_net_1\, Y => \address_7[28]\);
    
    \address_RNO[11]\ : MX2
      port map(A => N_20_0_i_0, B => addr_data_f2(11), S => 
        \state_0[0]_net_1\, Y => \address_7[11]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_21\ : AO1C
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, C => N_30_0, Y => N_32);
    
    \FSM_SELECT_ADDRESS.state7_0_I_73\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => state7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_35\ : XNOR2
      port map(A => \un2_nb_send_next[5]\, B => 
        nb_burst_available(5), Y => \DWACT_BL_EQUAL_0_E[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_2\ : XNOR2
      port map(A => \un2_nb_send_next[6]\, B => 
        nb_burst_available(6), Y => \DWACT_BL_EQUAL_0_E_0[0]\);
    
    un1_address_m38 : AX1
      port map(A => N_37_0, B => \addr_data_vector[86]\, C => 
        \addr_data_vector[87]\, Y => \un1_address[23]\);
    
    un1_address_m12 : AO13
      port map(A => N_5_0, B => address_0_sqmuxa, C => 
        \addr_data_vector[70]\, Y => N_13_0);
    
    un1_address_m59 : XNOR2
      port map(A => N_41, B => \addr_data_vector[88]\, Y => 
        \un1_address[24]\);
    
    \update_r[0]\ : DFN1P0
      port map(D => update_and_sel_3(4), CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \update_r_i[0]\);
    
    un2_nb_send_next_I_5 : XOR2
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        Y => \un2_nb_send_next[1]\);
    
    \address_RNO[17]\ : MX2
      port map(A => N_30_0_i_0, B => addr_data_f2(17), S => 
        \state_0[0]_net_1\, Y => \address_7[17]\);
    
    \address_RNO[5]\ : MX2
      port map(A => N_52_i_0, B => addr_data_f2(5), S => 
        \state_0[0]_net_1\, Y => \address_7[5]\);
    
    un1_address_m15 : OR3B
      port map(A => \addr_data_vector[71]\, B => 
        \addr_data_vector[72]\, C => N_13_0, Y => N_16_0);
    
    un1_address_m58 : XNOR2
      port map(A => N_37_0, B => \addr_data_vector[86]\, Y => 
        \un1_address[22]\);
    
    un2_nb_send_next_I_56 : XOR2
      port map(A => N_4, B => \nb_send[10]_net_1\, Y => 
        \un2_nb_send_next[10]\);
    
    \address_RNID894[14]\ : MX2C
      port map(A => addr_data_vector_11, B => 
        \addr_data_vector[78]\, S => sel_data_1(1), Y => N_1321);
    
    un2_nb_send_next_I_41 : AND2
      port map(A => \nb_send[6]_net_1\, B => \nb_send[7]_net_1\, 
        Y => \DWACT_FINC_E[3]\);
    
    un1_address_m41_m6_0_a2_6 : NOR3C
      port map(A => \addr_data_vector[86]\, B => 
        \addr_data_vector[85]\, C => m41_m6_0_a2_4, Y => 
        m41_m6_0_a2_6);
    
    \address_RNO[3]\ : MX2
      port map(A => N_50_i_0, B => addr_data_f2(3), S => 
        \state_0[0]_net_1\, Y => \address_7[3]\);
    
    \address[3]\ : DFN1C0
      port map(D => \address_7[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[67]\);
    
    un2_nb_send_next_I_34 : AND3
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        C => \nb_send[5]_net_1\, Y => \DWACT_FINC_E[2]\);
    
    un1_address_m64 : AX1C
      port map(A => \addr_data_vector[92]\, B => N_45, C => 
        \addr_data_vector[93]\, Y => \un1_address[29]\);
    
    \address_RNI58OA[9]\ : MX2C
      port map(A => addr_data_vector_6, B => 
        \addr_data_vector[73]\, S => sel_data_1(1), Y => N_1316);
    
    un1_address_m34 : XNOR2
      port map(A => N_34_0, B => \addr_data_vector[84]\, Y => 
        \un1_address[20]\);
    
    \address_RNO[30]\ : MX2
      port map(A => \un1_address[30]\, B => addr_data_f2(30), S
         => \state[0]_net_1\, Y => \address_7[30]\);
    
    un1_address_m26_m6_0_a2_2 : NOR2B
      port map(A => \addr_data_vector[74]\, B => 
        \addr_data_vector[75]\, Y => m26_m6_0_a2_2);
    
    \state_RNO_0[1]\ : OR2
      port map(A => status_full_ack(2), B => N_131, Y => 
        \state_ns_i_0[3]\);
    
    \nb_send[3]\ : DFN1E0C0
      port map(D => \nb_send_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[3]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_20\ : OR2A
      port map(A => nb_burst_available(10), B => 
        \un2_nb_send_next[10]\, Y => N_31);
    
    un1_address_m54 : XNOR2
      port map(A => N_23_0, B => \addr_data_vector[77]\, Y => 
        N_55_0_i_0);
    
    un1_address_m22 : OR3B
      port map(A => \addr_data_vector[75]\, B => 
        \addr_data_vector[76]\, C => N_19_0, Y => N_23_0);
    
    \address[7]\ : DFN1C0
      port map(D => \address_7[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[71]\);
    
    un2_nb_send_next_I_38 : XOR2
      port map(A => N_17, B => \nb_send[7]_net_1\, Y => 
        \un2_nb_send_next[7]\);
    
    \nb_send[5]\ : DFN1E0C0
      port map(D => \nb_send_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[5]_net_1\);
    
    \nb_send_RNO[5]\ : NOR2B
      port map(A => \un2_nb_send_next[5]\, B => state7, Y => 
        \nb_send_5[5]\);
    
    \address_RNIF894[15]\ : MX2C
      port map(A => addr_data_vector_12, B => 
        \addr_data_vector[79]\, S => sel_data_1(1), Y => N_1322);
    
    un1_address_m25 : XNOR2
      port map(A => N_25_0, B => \addr_data_vector[79]\, Y => 
        N_26_0_i_0);
    
    \state[3]\ : DFN1C0
      port map(D => N_113, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[3]_net_1\);
    
    \update_r_RNI3KV4[0]\ : OR2B
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => un3_update_r);
    
    \update_r[1]\ : DFN1C0
      port map(D => update_and_sel_3(5), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \update_r[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_17\ : OR2A
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, Y => N_28);
    
    \FSM_SELECT_ADDRESS.state7_0_I_43\ : AO1A
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => nb_burst_available(5), Y => 
        \ACT_LT2_E[2]\);
    
    \update_r_RNI3KV4_0[0]\ : OR2
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => \un1_state_12_3_0[4]\);
    
    un1_address_m40 : OR3B
      port map(A => \addr_data_vector[86]\, B => 
        \addr_data_vector[87]\, C => N_37_0, Y => N_41);
    
    \address_RNIIO94[31]\ : MX2C
      port map(A => addr_data_vector_28, B => 
        \addr_data_vector[95]\, S => sel_data_0(1), Y => N_1296);
    
    un1_address_m57 : AX1
      port map(A => N_34_0, B => \addr_data_vector[84]\, C => 
        \addr_data_vector[85]\, Y => \un1_address[21]\);
    
    un2_nb_send_next_I_8 : NOR2B
      port map(A => \nb_send[1]_net_1\, B => \nb_send[0]_net_1\, 
        Y => N_38);
    
    \FSM_SELECT_ADDRESS.state7_0_I_23\ : AO1C
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), C => N_28, Y => N_34);
    
    \FSM_SELECT_ADDRESS.state7_0_I_26\ : OA1A
      port map(A => N_32, B => N_34, C => N_33, Y => N_37);
    
    \address_RNO[22]\ : MX2
      port map(A => \un1_address[22]\, B => addr_data_f2(22), S
         => \state[0]_net_1\, Y => \address_7[22]\);
    
    un2_nb_send_next_I_27 : AND2
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        Y => \DWACT_FINC_E[1]\);
    
    un1_address_m49 : AX1C
      port map(A => \addr_data_vector[66]\, B => 
        \un1_state_12[4]\, C => \addr_data_vector[67]\, Y => 
        N_50_i_0);
    
    \address[9]\ : DFN1C0
      port map(D => \address_7[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[73]\);
    
    \address_RNO[18]\ : MX2
      port map(A => \un1_address[18]\, B => addr_data_f2(18), S
         => \state_0[0]_net_1\, Y => \address_7[18]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \address_RNO[7]\ : MX2
      port map(A => N_1_i_0, B => addr_data_f2(7), S => 
        \state_0[0]_net_1\, Y => \address_7[7]\);
    
    un1_address_m48 : AX1C
      port map(A => \addr_data_vector[94]\, B => N_47, C => 
        \addr_data_vector[95]\, Y => N_49_i_0);
    
    \address[6]\ : DFN1C0
      port map(D => \address_7[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[70]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_59\ : OR2A
      port map(A => \un2_nb_send_next[3]\, B => 
        nb_burst_available(3), Y => \ACT_LT4_E[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_1\ : XNOR2
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => \DWACT_BL_EQUAL_0_E[4]\);
    
    status_full_err_RNO : OR3
      port map(A => \state[3]_net_1\, B => \state[4]_net_1\, C
         => N_130, Y => N_110);
    
    \state_0[0]\ : DFN1C0
      port map(D => N_118, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state_0[0]_net_1\);
    
    \address_RNO[8]\ : MX2
      port map(A => N_15_0_i_0, B => addr_data_f2(8), S => 
        \state_0[0]_net_1\, Y => \address_7[8]\);
    
    un1_address_m36 : OR3B
      port map(A => \addr_data_vector[84]\, B => 
        \addr_data_vector[85]\, C => N_34_0, Y => N_37_0);
    
    un2_nb_send_next_I_52 : XOR2
      port map(A => N_7, B => \nb_send[9]_net_1\, Y => 
        \un2_nb_send_next[9]\);
    
    \address[11]\ : DFN1C0
      port map(D => \address_7[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[75]\);
    
    \state_RNIHABE[1]\ : NOR2A
      port map(A => status_full_ack(2), B => N_131, Y => N_118);
    
    \address[31]\ : DFN1C0
      port map(D => \address_7[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[95]\);
    
    \state_RNISHSP8[3]\ : OR2B
      port map(A => \state[3]_net_1\, B => state7, Y => 
        \un1_state_12_2[4]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_55\ : OR2A
      port map(A => nb_burst_available(2), B => 
        \un2_nb_send_next[2]\, Y => \ACT_LT4_E[4]\);
    
    un1_address_m56 : XNOR2
      port map(A => N_31_0, B => \addr_data_vector[82]\, Y => 
        \un1_address[18]\);
    
    \address_RNO[2]\ : MX2
      port map(A => N_40_i_0, B => addr_data_f2(2), S => 
        \state_0[0]_net_1\, Y => \address_7[2]\);
    
    un1_address_m44 : NOR3C
      port map(A => \addr_data_vector[90]\, B => N_43, C => 
        \addr_data_vector[91]\, Y => N_45);
    
    \address_RNO[4]\ : MX2
      port map(A => N_51_i_0, B => addr_data_f2(4), S => 
        \state_0[0]_net_1\, Y => \address_7[4]\);
    
    un2_nb_send_next_I_19 : NOR2B
      port map(A => \nb_send[3]_net_1\, B => \DWACT_FINC_E[0]\, Y
         => N_30);
    
    \address_RNO[25]\ : MX2
      port map(A => \un1_address[25]\, B => addr_data_f2(25), S
         => \state[0]_net_1\, Y => \address_7[25]\);
    
    \address[21]\ : DFN1C0
      port map(D => \address_7[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[85]\);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    un1_address_m62 : AX1C
      port map(A => \addr_data_vector[90]\, B => N_43, C => 
        \addr_data_vector[91]\, Y => \un1_address[27]\);
    
    un1_address_m32 : AX1
      port map(A => N_31_0, B => \addr_data_vector[82]\, C => 
        \addr_data_vector[83]\, Y => \un1_address[19]\);
    
    un1_address_m12_e : OR3C
      port map(A => \addr_data_vector[68]\, B => N_69, C => 
        \addr_data_vector[69]\, Y => N_5_0);
    
    un2_nb_send_next_I_9 : XOR2
      port map(A => N_38, B => \nb_send[2]_net_1\, Y => 
        \un2_nb_send_next[2]\);
    
    \state[1]\ : DFN1C0
      port map(D => N_116, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[1]_net_1\);
    
    \address[17]\ : DFN1C0
      port map(D => \address_7[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[81]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_52\ : OR2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[1]\);
    
    un1_address_m65 : XOR2
      port map(A => N_47, B => \addr_data_vector[94]\, Y => 
        \un1_address[30]\);
    
    un1_address_m52 : XNOR2
      port map(A => N_13_0, B => \addr_data_vector[71]\, Y => 
        N_1_i_0);
    
    \address[27]\ : DFN1C0
      port map(D => \address_7[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[91]\);
    
    \state_RNO[3]\ : NOR2A
      port map(A => \state[4]_net_1\, B => N_129, Y => N_113);
    
    un1_address_m21 : AX1
      port map(A => N_19_0, B => \addr_data_vector[75]\, C => 
        \addr_data_vector[76]\, Y => N_22_0_i_0);
    
    \nb_send_RNO[4]\ : NOR2B
      port map(A => \un2_nb_send_next[4]\, B => state7, Y => 
        \nb_send_5[4]\);
    
    \nb_send_RNO[10]\ : NOR2B
      port map(A => \un2_nb_send_next[10]\, B => state7, Y => 
        \nb_send_5[10]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_18\ : OR2A
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => N_29);
    
    un1_address_m55 : AX1
      port map(A => N_23_0, B => \addr_data_vector[77]\, C => 
        \addr_data_vector[78]\, Y => N_56_0_i_0);
    
    \address_RNO[31]\ : MX2
      port map(A => N_49_i_0, B => addr_data_f2(31), S => 
        \state[0]_net_1\, Y => \address_7[31]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_61\ : AOI1A
      port map(A => \ACT_LT4_E[3]\, B => \ACT_LT4_E[6]\, C => 
        \ACT_LT4_E[10]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\);
    
    un1_address_m10_e : NOR3C
      port map(A => \addr_data_vector[66]\, B => 
        \un1_state_12[4]\, C => \addr_data_vector[67]\, Y => N_69);
    
    \FSM_SELECT_ADDRESS.state7_0_I_34\ : XNOR2
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), Y => \DWACT_BL_EQUAL_0_E[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_6\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E_0[0]\, B => 
        \DWACT_BL_EQUAL_0_E_0[1]\, C => \DWACT_BL_EQUAL_0_E[2]\, 
        Y => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\);
    
    \address_RNO[12]\ : MX2
      port map(A => N_22_0_i_0, B => addr_data_f2(12), S => 
        \state_0[0]_net_1\, Y => \address_7[12]\);
    
    un2_nb_send_next_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \nb_send[6]_net_1\, Y => N_17);
    
    un2_nb_send_next_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_12);
    
    \FSM_SELECT_ADDRESS.state7_0_I_3\ : XNOR2
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => \DWACT_BL_EQUAL_0_E[2]\);
    
    status_full_RNO : OR2
      port map(A => \state[2]_net_1\, B => N_126, Y => 
        un1_state_11);
    
    \address[1]\ : DFN1E1C0
      port map(D => addr_data_f2(1), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        addr_data_vector_62);
    
    \status_full\ : DFN1E1C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_11, Q => status_full(2));
    
    un1_address_m63 : XOR2
      port map(A => N_45, B => \addr_data_vector[92]\, Y => 
        \un1_address[28]\);
    
    un1_address_m33 : OR3B
      port map(A => \addr_data_vector[82]\, B => 
        \addr_data_vector[83]\, C => N_31_0, Y => N_34_0);
    
    un1_address_m26_m6_0_a2_4 : NOR3C
      port map(A => \addr_data_vector[71]\, B => 
        \addr_data_vector[79]\, C => \addr_data_vector[78]\, Y
         => m26_m6_0_a2_4);
    
    un2_nb_send_next_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    un1_address_m41_m6_0_a2_2 : NOR2B
      port map(A => \addr_data_vector[83]\, B => 
        \addr_data_vector[84]\, Y => m41_m6_0_a2_2);
    
    un1_address_m41_m6_0_a2_1 : NOR2B
      port map(A => \addr_data_vector[81]\, B => 
        \addr_data_vector[82]\, Y => m41_m6_0_a2_1);
    
    \address_RNO[20]\ : MX2
      port map(A => \un1_address[20]\, B => addr_data_f2(20), S
         => \state[0]_net_1\, Y => \address_7[20]\);
    
    un1_address_m46 : NOR3C
      port map(A => \addr_data_vector[92]\, B => N_45, C => 
        \addr_data_vector[93]\, Y => N_47);
    
    \nb_send[8]\ : DFN1E0C0
      port map(D => \nb_send_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[8]_net_1\);
    
    un1_address_m53 : AX1
      port map(A => N_16_0, B => \addr_data_vector[73]\, C => 
        \addr_data_vector[74]\, Y => N_54_0_i_0);
    
    \state_RNIVJCD[1]\ : NOR2
      port map(A => \state[2]_net_1\, B => \state[1]_net_1\, Y
         => N_131);
    
    \nb_send[1]\ : DFN1E0C0
      port map(D => \nb_send_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_60\ : AOI1A
      port map(A => \ACT_LT4_E[7]\, B => \ACT_LT4_E[8]\, C => 
        \ACT_LT4_E[5]\, Y => \ACT_LT4_E[10]\);
    
    un1_address_m41_m6_0_a2_4 : NOR3C
      port map(A => \addr_data_vector[80]\, B => 
        \addr_data_vector[88]\, C => \addr_data_vector[87]\, Y
         => m41_m6_0_a2_4);
    
    \state_RNIH9F11[2]\ : NOR2B
      port map(A => \state[2]_net_1\, B => N_129, Y => N_130);
    
    \state_RNO_1[4]\ : OR3A
      port map(A => \state_0[0]_net_1\, B => \state[3]_net_1\, C
         => \state[2]_net_1\, Y => N_124);
    
    \address_RNO[15]\ : MX2
      port map(A => N_26_0_i_0, B => addr_data_f2(15), S => 
        \state_0[0]_net_1\, Y => \address_7[15]\);
    
    un2_nb_send_next_I_20 : XOR2
      port map(A => N_30, B => \nb_send[4]_net_1\, Y => 
        \un2_nb_send_next[4]\);
    
    un1_address_m42 : NOR3B
      port map(A => m41_m6_0_a2_7, B => \addr_data_vector[89]\, C
         => N_27_0_i_0, Y => N_43);
    
    \FSM_SELECT_ADDRESS.state7_0_I_68\ : AO1
      port map(A => \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, B => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, C => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, Y => 
        \DWACT_COMP0_E[2]\);
    
    \address_RNIVHIB[8]\ : MX2C
      port map(A => addr_data_vector_5, B => 
        \addr_data_vector[72]\, S => sel_data(1), Y => N_1329);
    
    un2_nb_send_next_I_16 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\ is

    port( nb_burst_available  : in    std_logic_vector(10 downto 0);
          status_full_err     : out   std_logic_vector(0 to 0);
          status_full         : out   std_logic_vector(0 to 0);
          sel_data            : in    std_logic_vector(1 to 1);
          sel_data_1          : in    std_logic_vector(1 to 1);
          sel_data_0          : in    std_logic_vector(1 to 1);
          update_and_sel_7    : in    std_logic_vector(1 downto 0);
          addr_data_f0        : in    std_logic_vector(31 downto 0);
          status_full_ack     : in    std_logic_vector(0 to 0);
          addr_data_vector_69 : in    std_logic;
          addr_data_vector_68 : in    std_logic;
          addr_data_vector_66 : in    std_logic;
          addr_data_vector_77 : in    std_logic;
          addr_data_vector_75 : in    std_logic;
          addr_data_vector_86 : in    std_logic;
          addr_data_vector_85 : in    std_logic;
          addr_data_vector_84 : in    std_logic;
          addr_data_vector_83 : in    std_logic;
          addr_data_vector_82 : in    std_logic;
          addr_data_vector_81 : in    std_logic;
          addr_data_vector_80 : in    std_logic;
          addr_data_vector_92 : in    std_logic;
          addr_data_vector_90 : in    std_logic;
          addr_data_vector_88 : in    std_logic;
          addr_data_vector_87 : in    std_logic;
          addr_data_vector_94 : in    std_logic;
          addr_data_vector_65 : in    std_logic;
          addr_data_vector_64 : in    std_logic;
          addr_data_vector_3  : out   std_logic;
          addr_data_vector_31 : out   std_logic;
          addr_data_vector_14 : out   std_logic;
          addr_data_vector_15 : out   std_logic;
          addr_data_vector_27 : out   std_logic;
          addr_data_vector_29 : out   std_logic;
          addr_data_vector_25 : out   std_logic;
          addr_data_vector_6  : out   std_logic;
          addr_data_vector_8  : out   std_logic;
          addr_data_vector_7  : out   std_logic;
          addr_data_vector_10 : out   std_logic;
          addr_data_vector_9  : out   std_logic;
          addr_data_vector_12 : out   std_logic;
          N_1326              : out   std_logic;
          N_1325              : out   std_logic;
          N_1323              : out   std_logic;
          N_1320              : out   std_logic;
          N_1318              : out   std_logic;
          N_1315              : out   std_logic;
          N_1314              : out   std_logic;
          N_1313              : out   std_logic;
          N_1312              : out   std_logic;
          N_1311              : out   std_logic;
          N_1310              : out   std_logic;
          N_1309              : out   std_logic;
          N_1307              : out   std_logic;
          N_1305              : out   std_logic;
          N_1303              : out   std_logic;
          N_1302              : out   std_logic;
          N_1295              : out   std_logic;
          N_1280              : out   std_logic;
          N_1279              : out   std_logic;
          HRESETn_c           : in    std_logic;
          HCLK_c              : in    std_logic
        );

end 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\ is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \state_0[0]_net_1\, \state_RNIBABE[1]_net_1\, N_38, 
        \nb_send[1]_net_1\, \nb_send[0]_net_1\, N_30, 
        \nb_send[3]_net_1\, \DWACT_FINC_E[0]\, N_7, 
        \nb_send[8]_net_1\, \DWACT_FINC_E[4]\, m40_m6_0_a2_7, 
        m40_m6_0_a2_6, m37_m6_0_a2_4_i, m40_m6_0_a2_3, 
        m40_m6_0_a2_2, m40_m6_0_a2_4, \addr_data_vector[13]\, 
        \addr_data_vector[23]\, m40_m6_0_a2_1, 
        \addr_data_vector[11]\, m23_m7_i_5, m23_m7_i_2, 
        m23_m7_i_1, m23_m7_i_3, \addr_data_vector[7]\, 
        \addr_data_vector[12]\, \addr_data_vector[10]\, 
        \addr_data_vector[8]\, \addr_data_vector[9]\, 
        ADD_32x32_fast_I164_Y_0_0, address_0_sqmuxa, 
        \un1_state_12_3_0[4]\, \update_r_i[0]\, 
        \update_r[1]_net_1\, address_0_sqmuxa_0, \state[3]_net_1\, 
        un3_update_r, un1_state_5_i_0, \state[4]_net_1\, 
        \state_ns_i_0[3]\, N_85, address_7_31_m6_e_3, 
        \addr_data_vector[30]\, address_7_31_m6_e_1, 
        address_7_31_m6_e_2, \addr_data_vector[28]\, 
        \addr_data_vector[26]\, m37_m6_0_a2_4_6, 
        \addr_data_vector[20]\, \addr_data_vector[19]\, 
        m37_m6_0_a2_4_4, m37_m6_0_a2_4_5, \addr_data_vector[16]\, 
        m37_m6_0_a2_4_2, \addr_data_vector[22]\, 
        \addr_data_vector[21]\, \addr_data_vector[17]\, 
        \addr_data_vector[18]\, \un1_address[6]\, N_5_0, 
        \state_RNO_0[1]_net_1\, N_83_i, \state[1]_net_1\, 
        \state_ns[0]\, N_79, N_78, \un1_state_12_2[4]\, N_64, 
        N_84, \state[2]_net_1\, state7, \address_RNO_2_0[31]\, 
        m23_m7_i, m23_N_10, m23_m7_i_a5, \addr_data_vector[6]\, 
        \address_7[31]\, \address_RNO_0_0[31]\, 
        \address_RNO_1_0[31]\, N_42, \addr_data_vector[31]\, N_2, 
        \addr_data_vector[2]\, N_4_0, \addr_data_vector[4]\, 
        N_15_0_i_0, N_13_0, N_16_0, N_17_0_i_0, N_19_0, 
        N_20_0_i_0, N_21_0, N_22_0_i_0, N_26_0_i_0, 
        \addr_data_vector[14]\, \addr_data_vector[15]\, N_27_0, 
        N_28_0_i_0, N_30_0_i_0, N_31_0, \un1_address[19]\, N_34_0, 
        \un1_address[20]\, N_36_0, \un1_address[23]\, N_40_i_0, 
        \addr_data_vector[24]\, N_44, \addr_data_vector[25]\, 
        N_46, \addr_data_vector[27]\, N_50_i_0, 
        \addr_data_vector[3]\, N_51_i_0, N_52_i_0, 
        \addr_data_vector[5]\, N_1_i_0, N_54_0_i_0, N_55_0_i_0, 
        \un1_address[18]\, \un1_address[21]\, \un1_address[22]\, 
        \un1_address[24]\, \un1_address[25]\, \un1_address[26]\, 
        \un1_address[27]\, \un1_address[28]\, \un1_address[29]\, 
        \addr_data_vector[29]\, \un1_address[30]\, \address_7[2]\, 
        \address_7[3]\, \address_7[4]\, \address_7[5]\, 
        \address_7[6]\, \address_7[7]\, \address_7[8]\, 
        \address_7[9]\, \address_7[10]\, \address_7[11]\, 
        \address_7[12]\, \address_7[13]\, \address_7[15]\, 
        \address_7[16]\, \address_7[17]\, \state[0]_net_1\, 
        \address_7[18]\, \address_7[19]\, \address_7[20]\, 
        \address_7[21]\, \address_7[22]\, \address_7[23]\, 
        \address_7[24]\, \address_7[25]\, \address_7[26]\, 
        \address_7[27]\, \address_7[28]\, \address_7[29]\, 
        \address_7[30]\, N_56_0_i_0, un1_state_9, \nb_send_5[0]\, 
        \nb_send_5[1]\, \un2_nb_send_next[1]\, \nb_send_5[2]\, 
        \un2_nb_send_next[2]\, \nb_send_5[3]\, 
        \un2_nb_send_next[3]\, \nb_send_5[4]\, 
        \un2_nb_send_next[4]\, \nb_send_5[5]\, 
        \un2_nb_send_next[5]\, \nb_send_5[6]\, 
        \un2_nb_send_next[6]\, \nb_send_5[7]\, 
        \un2_nb_send_next[7]\, \nb_send_5[8]\, 
        \un2_nb_send_next[8]\, \nb_send_5[9]\, 
        \un2_nb_send_next[9]\, \nb_send_5[10]\, 
        \un2_nb_send_next[10]\, N_80, \state_RNO_1[3]\, 
        \state_ns[2]\, un1_state_11, \address_7[14]\, 
        \addr_data_vector[0]\, \addr_data_vector[1]\, 
        \nb_send[2]_net_1\, \nb_send[4]_net_1\, 
        \nb_send[5]_net_1\, \nb_send[6]_net_1\, 
        \nb_send[7]_net_1\, \nb_send[9]_net_1\, 
        \nb_send[10]_net_1\, N_4, \DWACT_FINC_E[2]\, 
        \DWACT_FINC_E[3]\, N_12, N_17, N_22, \DWACT_FINC_E[1]\, 
        N_27, N_35, \DWACT_COMP0_E[1]\, \DWACT_COMP0_E[2]\, 
        \DWACT_COMP0_E[0]\, \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, \ACT_LT4_E[3]\, 
        \ACT_LT4_E[6]\, \ACT_LT4_E[10]\, \ACT_LT4_E[7]\, 
        \ACT_LT4_E[8]\, \ACT_LT4_E[5]\, \ACT_LT4_E[4]\, 
        \ACT_LT4_E[0]\, \ACT_LT4_E[1]\, \ACT_LT4_E[2]\, 
        \ACT_LT2_E[0]\, \ACT_LT2_E[1]\, \ACT_LT2_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, N_37, 
        N_36, N_35_0, N_32, N_34, N_33, N_31, N_28, N_29, N_30_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, 
        \DWACT_BL_EQUAL_0_E[4]\, \DWACT_BL_EQUAL_0_E[3]\, 
        \DWACT_BL_EQUAL_0_E_0[0]\, \DWACT_BL_EQUAL_0_E_0[1]\, 
        \DWACT_BL_EQUAL_0_E[2]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    addr_data_vector_3 <= \addr_data_vector[3]\;
    addr_data_vector_31 <= \addr_data_vector[31]\;
    addr_data_vector_14 <= \addr_data_vector[14]\;
    addr_data_vector_15 <= \addr_data_vector[15]\;
    addr_data_vector_27 <= \addr_data_vector[27]\;
    addr_data_vector_29 <= \addr_data_vector[29]\;
    addr_data_vector_25 <= \addr_data_vector[25]\;
    addr_data_vector_6 <= \addr_data_vector[6]\;
    addr_data_vector_8 <= \addr_data_vector[8]\;
    addr_data_vector_7 <= \addr_data_vector[7]\;
    addr_data_vector_10 <= \addr_data_vector[10]\;
    addr_data_vector_9 <= \addr_data_vector[9]\;
    addr_data_vector_12 <= \addr_data_vector[12]\;

    \address[16]\ : DFN1C0
      port map(D => \address_7[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[16]\);
    
    \address[10]\ : DFN1C0
      port map(D => \address_7[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[10]\);
    
    \state[0]\ : DFN1C0
      port map(D => \state_RNIBABE[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state[0]_net_1\);
    
    \address[30]\ : DFN1C0
      port map(D => \address_7[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[30]\);
    
    un1_address_m45 : NOR3C
      port map(A => \addr_data_vector[27]\, B => N_44, C => 
        \addr_data_vector[28]\, Y => N_46);
    
    \address_RNO[26]\ : MX2
      port map(A => \un1_address[26]\, B => addr_data_f0(26), S
         => \state[0]_net_1\, Y => \address_7[26]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_25\ : AO1C
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_31, Y => N_36);
    
    un1_address_m61 : AX1C
      port map(A => \addr_data_vector[25]\, B => N_42, C => 
        \addr_data_vector[26]\, Y => \un1_address[26]\);
    
    \address_RNIN894[19]\ : MX2C
      port map(A => \addr_data_vector[19]\, B => 
        addr_data_vector_83, S => sel_data_1(1), Y => N_1312);
    
    un1_address_m37_m6_0_a2_4_6 : NOR3C
      port map(A => \addr_data_vector[20]\, B => 
        \addr_data_vector[19]\, C => m37_m6_0_a2_4_4, Y => 
        m37_m6_0_a2_4_6);
    
    un1_address_m37_m6_0_a2_4 : OR2B
      port map(A => m37_m6_0_a2_4_6, B => m37_m6_0_a2_4_5, Y => 
        m37_m6_0_a2_4_i);
    
    \address[26]\ : DFN1C0
      port map(D => \address_7[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[26]\);
    
    \address[20]\ : DFN1C0
      port map(D => \address_7[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[20]\);
    
    \address_RNIK7MA[1]\ : MX2C
      port map(A => \addr_data_vector[1]\, B => 
        addr_data_vector_65, S => sel_data_0(1), Y => N_1280);
    
    \state_RNI9QRU8_0[3]\ : OR2B
      port map(A => address_0_sqmuxa_0, B => state7, Y => 
        address_0_sqmuxa);
    
    \FSM_SELECT_ADDRESS.state7_0_I_42\ : AO1C
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => \un2_nb_send_next[5]\, Y => 
        \ACT_LT2_E[1]\);
    
    \address_RNIPPHB[5]\ : MX2C
      port map(A => \addr_data_vector[5]\, B => 
        addr_data_vector_69, S => sel_data(1), Y => N_1326);
    
    \FSM_SELECT_ADDRESS.state7_0_I_57\ : NOR2A
      port map(A => \ACT_LT4_E[4]\, B => \ACT_LT4_E[5]\, Y => 
        \ACT_LT4_E[6]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_36\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[1]\, B => 
        \DWACT_BL_EQUAL_0_E[0]\, Y => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\);
    
    un1_address_m51 : XOR2
      port map(A => N_4_0, B => \addr_data_vector[5]\, Y => 
        N_52_i_0);
    
    \address[12]\ : DFN1C0
      port map(D => \address_7[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[12]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_22\ : OA1A
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_29, Y => N_33);
    
    \address_RNO[29]\ : MX2
      port map(A => \un1_address[29]\, B => addr_data_f0(29), S
         => \state[0]_net_1\, Y => \address_7[29]\);
    
    \update_r_RNIVJV4[0]\ : OR2B
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => un3_update_r);
    
    \FSM_SELECT_ADDRESS.state7_0_I_8\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, B => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, Y => 
        \DWACT_COMP0_E[1]\);
    
    un1_address_m19 : XNOR2
      port map(A => N_19_0, B => \addr_data_vector[11]\, Y => 
        N_20_0_i_0);
    
    \address[22]\ : DFN1C0
      port map(D => \address_7[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[22]\);
    
    \address_RNO[23]\ : MX2
      port map(A => \un1_address[23]\, B => addr_data_f0(23), S
         => \state[0]_net_1\, Y => \address_7[23]\);
    
    \address[2]\ : DFN1C0
      port map(D => \address_7[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[2]\);
    
    un2_nb_send_next_I_13 : XOR2
      port map(A => N_35, B => \nb_send[3]_net_1\, Y => 
        \un2_nb_send_next[3]\);
    
    un1_address_m43 : NOR3C
      port map(A => \addr_data_vector[25]\, B => N_42, C => 
        \addr_data_vector[26]\, Y => N_44);
    
    \FSM_SELECT_ADDRESS.state7_0_I_54\ : AOI1A
      port map(A => \ACT_LT4_E[0]\, B => \ACT_LT4_E[1]\, C => 
        \ACT_LT4_E[2]\, Y => \ACT_LT4_E[3]\);
    
    \address_RNO[24]\ : MX2
      port map(A => \un1_address[24]\, B => addr_data_f0(24), S
         => \state[0]_net_1\, Y => \address_7[24]\);
    
    \address_RNO[10]\ : MX2
      port map(A => N_54_0_i_0, B => addr_data_f0(10), S => 
        \state_0[0]_net_1\, Y => \address_7[10]\);
    
    \status_full_err\ : DFN1E0C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_64, Q => status_full_err(0));
    
    un2_nb_send_next_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \nb_send[8]_net_1\, C
         => \nb_send[9]_net_1\, Y => N_4);
    
    un1_address_m18 : OR3B
      port map(A => \addr_data_vector[9]\, B => 
        \addr_data_vector[10]\, C => N_16_0, Y => N_19_0);
    
    \nb_send_RNO[1]\ : NOR2B
      port map(A => \un2_nb_send_next[1]\, B => state7, Y => 
        \nb_send_5[1]\);
    
    \state_RNIF9F11[2]\ : NOR2A
      port map(A => \state[2]_net_1\, B => N_83_i, Y => N_84);
    
    un1_address_ADD_32x32_fast_I164_Y_0_0 : XNOR2
      port map(A => \addr_data_vector[6]\, B => address_0_sqmuxa, 
        Y => ADD_32x32_fast_I164_Y_0_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_51\ : NOR2B
      port map(A => \nb_send[0]_net_1\, B => 
        nb_burst_available(0), Y => \ACT_LT4_E[0]\);
    
    un2_nb_send_next_I_31 : XOR2
      port map(A => N_22, B => \nb_send[6]_net_1\, Y => 
        \un2_nb_send_next[6]\);
    
    \nb_send[9]\ : DFN1E0C0
      port map(D => \nb_send_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[9]_net_1\);
    
    \address_RNO[9]\ : MX2
      port map(A => N_17_0_i_0, B => addr_data_f0(9), S => 
        \state_0[0]_net_1\, Y => \address_7[9]\);
    
    \address[5]\ : DFN1C0
      port map(D => \address_7[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[5]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_5\ : XNOR2
      port map(A => \un2_nb_send_next[7]\, B => 
        nb_burst_available(7), Y => \DWACT_BL_EQUAL_0_E_0[1]\);
    
    \address[15]\ : DFN1C0
      port map(D => \address_7[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[15]\);
    
    \address[13]\ : DFN1C0
      port map(D => \address_7[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[13]\);
    
    un1_address_m20 : NOR2A
      port map(A => \addr_data_vector[11]\, B => N_19_0, Y => 
        N_21_0);
    
    \state[4]\ : DFN1P0
      port map(D => \state_ns[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[4]_net_1\);
    
    \address_RNIJ894[17]\ : MX2C
      port map(A => \addr_data_vector[17]\, B => 
        addr_data_vector_81, S => sel_data_1(1), Y => N_1310);
    
    \nb_send_RNO[9]\ : NOR2B
      port map(A => \un2_nb_send_next[9]\, B => state7, Y => 
        \nb_send_5[9]\);
    
    \address[19]\ : DFN1C0
      port map(D => \address_7[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[19]\);
    
    \address[25]\ : DFN1C0
      port map(D => \address_7[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[25]\);
    
    un2_nb_send_next_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => \nb_send[5]_net_1\, Y => N_22);
    
    \address[23]\ : DFN1C0
      port map(D => \address_7[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[23]\);
    
    un1_address_m14 : AX1
      port map(A => N_13_0, B => \addr_data_vector[7]\, C => 
        \addr_data_vector[8]\, Y => N_15_0_i_0);
    
    un1_address_m29 : AX1
      port map(A => N_27_0, B => \addr_data_vector[16]\, C => 
        \addr_data_vector[17]\, Y => N_30_0_i_0);
    
    un2_nb_send_next_I_12 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => N_35);
    
    \FSM_SELECT_ADDRESS.state7_0_I_19\ : NOR2A
      port map(A => nb_burst_available(6), B => 
        \un2_nb_send_next[6]\, Y => N_30_0);
    
    \address_RNO_2[31]\ : NOR3B
      port map(A => address_7_31_m6_e_3, B => address_7_31_m6_e_2, 
        C => \state_0[0]_net_1\, Y => \address_RNO_2_0[31]\);
    
    \address[29]\ : DFN1C0
      port map(D => \address_7[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[29]\);
    
    \address[18]\ : DFN1C0
      port map(D => \address_7[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[18]\);
    
    \nb_send_RNO[6]\ : NOR2B
      port map(A => \un2_nb_send_next[6]\, B => state7, Y => 
        \nb_send_5[6]\);
    
    \address_RNO[21]\ : MX2
      port map(A => \un1_address[21]\, B => addr_data_f0(21), S
         => \state[0]_net_1\, Y => \address_7[21]\);
    
    \address_RNO[16]\ : MX2
      port map(A => N_28_0_i_0, B => addr_data_f0(16), S => 
        \state_0[0]_net_1\, Y => \address_7[16]\);
    
    un2_nb_send_next_I_51 : NOR2B
      port map(A => \nb_send[8]_net_1\, B => \DWACT_FINC_E[4]\, Y
         => N_7);
    
    \address_RNIH894[16]\ : MX2C
      port map(A => \addr_data_vector[16]\, B => 
        addr_data_vector_80, S => sel_data_1(1), Y => N_1309);
    
    \address[0]\ : DFN1E1C0
      port map(D => addr_data_f0(0), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        \addr_data_vector[0]\);
    
    status_full_err_RNO_0 : OR2
      port map(A => \state[4]_net_1\, B => \state[3]_net_1\, Y
         => un1_state_5_i_0);
    
    \state_RNIRJCD[1]\ : NOR2
      port map(A => \state[2]_net_1\, B => \state[1]_net_1\, Y
         => N_85);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_address_m41 : NOR3B
      port map(A => m40_m6_0_a2_7, B => \addr_data_vector[24]\, C
         => N_13_0, Y => N_42);
    
    \address_RNO[27]\ : MX2
      port map(A => \un1_address[27]\, B => addr_data_f0(27), S
         => \state[0]_net_1\, Y => \address_7[27]\);
    
    \address[4]\ : DFN1C0
      port map(D => \address_7[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[4]\);
    
    \address[28]\ : DFN1C0
      port map(D => \address_7[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[28]\);
    
    un1_address_m1 : NOR3A
      port map(A => \addr_data_vector[2]\, B => 
        \un1_state_12_2[4]\, C => \un1_state_12_3_0[4]\, Y => N_2);
    
    \FSM_SELECT_ADDRESS.state7_0_I_7\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[4]\, B => 
        \DWACT_BL_EQUAL_0_E[3]\, Y => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\);
    
    \nb_send_RNO[2]\ : NOR2B
      port map(A => \un2_nb_send_next[2]\, B => state7, Y => 
        \nb_send_5[2]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \state_RNO_0[4]\ : OR3A
      port map(A => N_85, B => \state[3]_net_1\, C => N_83_i, Y
         => N_79);
    
    \address_RNO_1[31]\ : XNOR2
      port map(A => N_42, B => \addr_data_vector[31]\, Y => 
        \address_RNO_1_0[31]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_58\ : NOR2A
      port map(A => \un2_nb_send_next[2]\, B => 
        nb_burst_available(2), Y => \ACT_LT4_E[7]\);
    
    \nb_send_RNO[7]\ : NOR2B
      port map(A => \un2_nb_send_next[7]\, B => state7, Y => 
        \nb_send_5[7]\);
    
    un2_nb_send_next_I_24 : XOR2
      port map(A => N_27, B => \nb_send[5]_net_1\, Y => 
        \un2_nb_send_next[5]\);
    
    un2_nb_send_next_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \nb_send[3]_net_1\, C
         => \nb_send[4]_net_1\, Y => N_27);
    
    un1_address_ADD_32x32_fast_I164_Y_0 : XNOR2
      port map(A => ADD_32x32_fast_I164_Y_0_0, B => N_5_0, Y => 
        \un1_address[6]\);
    
    \address_RNO[19]\ : MX2
      port map(A => \un1_address[19]\, B => addr_data_f0(19), S
         => \state[0]_net_1\, Y => \address_7[19]\);
    
    \nb_send[7]\ : DFN1E0C0
      port map(D => \nb_send_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[7]_net_1\);
    
    \address_RNO[13]\ : MX2
      port map(A => N_55_0_i_0, B => addr_data_f0(13), S => 
        \state_0[0]_net_1\, Y => \address_7[13]\);
    
    \address[14]\ : DFN1C0
      port map(D => \address_7[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[14]\);
    
    un1_address_m23_m7_i_a5_0 : OR2B
      port map(A => N_5_0, B => address_0_sqmuxa, Y => m23_N_10);
    
    \state_RNO[1]\ : OA1B
      port map(A => N_83_i, B => \state[1]_net_1\, C => 
        \state_ns_i_0[3]\, Y => \state_RNO_0[1]_net_1\);
    
    \nb_send[0]\ : DFN1E0C0
      port map(D => \nb_send_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[0]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_53\ : AND2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[2]\);
    
    un1_address_m40_m6_0_a2_4 : NOR3C
      port map(A => \addr_data_vector[13]\, B => 
        \addr_data_vector[23]\, C => m40_m6_0_a2_1, Y => 
        m40_m6_0_a2_4);
    
    \nb_send[6]\ : DFN1E0C0
      port map(D => \nb_send_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[6]_net_1\);
    
    \nb_send[10]\ : DFN1E0C0
      port map(D => \nb_send_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[10]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_56\ : NOR2A
      port map(A => nb_burst_available(3), B => 
        \un2_nb_send_next[3]\, Y => \ACT_LT4_E[5]\);
    
    \address_RNO[14]\ : MX2
      port map(A => N_56_0_i_0, B => addr_data_f0(14), S => 
        \state[0]_net_1\, Y => \address_7[14]\);
    
    un1_address_m23_m7_i_a5 : AO1D
      port map(A => N_5_0, B => address_0_sqmuxa, C => 
        \addr_data_vector[6]\, Y => m23_m7_i_a5);
    
    \state_RNIA6SP8[3]\ : OR2B
      port map(A => \state[3]_net_1\, B => state7, Y => 
        \un1_state_12_2[4]\);
    
    \nb_send_RNO[3]\ : NOR2B
      port map(A => \un2_nb_send_next[3]\, B => state7, Y => 
        \nb_send_5[3]\);
    
    \nb_send[2]\ : DFN1E0C0
      port map(D => \nb_send_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[2]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_27\ : OA1
      port map(A => N_37, B => N_36, C => N_35_0, Y => 
        \DWACT_COMP0_E[0]\);
    
    \address[24]\ : DFN1C0
      port map(D => \address_7[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[24]\);
    
    un1_address_m27 : XNOR2
      port map(A => N_27_0, B => \addr_data_vector[16]\, Y => 
        N_28_0_i_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \address_RNO_0[31]\ : MX2C
      port map(A => \addr_data_vector[31]\, B => addr_data_f0(31), 
        S => \state_0[0]_net_1\, Y => \address_RNO_0_0[31]\);
    
    un1_address_m60 : XOR2
      port map(A => N_42, B => \addr_data_vector[25]\, Y => 
        \un1_address[25]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_44\ : AND3A
      port map(A => \ACT_LT2_E[0]\, B => \ACT_LT2_E[1]\, C => 
        \ACT_LT2_E[2]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\);
    
    un1_address_m30 : OR3B
      port map(A => \addr_data_vector[16]\, B => 
        \addr_data_vector[17]\, C => N_27_0, Y => N_31_0);
    
    \nb_send[4]\ : DFN1E0C0
      port map(D => \nb_send_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[4]_net_1\);
    
    un1_address_m16 : XNOR2
      port map(A => N_16_0, B => \addr_data_vector[9]\, Y => 
        N_17_0_i_0);
    
    un1_address_m37_m6_0_a2_4_2 : NOR2B
      port map(A => \addr_data_vector[17]\, B => 
        \addr_data_vector[18]\, Y => m37_m6_0_a2_4_2);
    
    un2_nb_send_next_I_45 : XOR2
      port map(A => N_12, B => \nb_send[8]_net_1\, Y => 
        \un2_nb_send_next[8]\);
    
    \nb_send_RNO[0]\ : NOR2A
      port map(A => state7, B => \nb_send[0]_net_1\, Y => 
        \nb_send_5[0]\);
    
    un1_address_m23_m7_i : OR3C
      port map(A => m23_N_10, B => m23_m7_i_5, C => m23_m7_i_a5, 
        Y => m23_m7_i);
    
    \state_RNI9QRU8[3]\ : AO1B
      port map(A => un3_update_r, B => state7, C => 
        \state[3]_net_1\, Y => un1_state_9);
    
    \nb_send_RNO[8]\ : NOR2B
      port map(A => \un2_nb_send_next[8]\, B => state7, Y => 
        \nb_send_5[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_41\ : AND2A
      port map(A => nb_burst_available(5), B => 
        \un2_nb_send_next[5]\, Y => \ACT_LT2_E[0]\);
    
    \state_RNO[4]\ : OR3C
      port map(A => N_79, B => N_78, C => \un1_state_12_2[4]\, Y
         => \state_ns[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_4\ : XNOR2
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), Y => \DWACT_BL_EQUAL_0_E[3]\);
    
    \address[8]\ : DFN1C0
      port map(D => \address_7[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[8]\);
    
    un1_address_m40_m6_0_a2_2 : NOR2B
      port map(A => \addr_data_vector[9]\, B => 
        \addr_data_vector[10]\, Y => m40_m6_0_a2_2);
    
    \address_RNIHG94[23]\ : MX2C
      port map(A => \addr_data_vector[23]\, B => 
        addr_data_vector_87, S => sel_data_1(1), Y => N_1302);
    
    un1_address_m50 : AX1C
      port map(A => \addr_data_vector[3]\, B => N_2, C => 
        \addr_data_vector[4]\, Y => N_51_i_0);
    
    un1_address_m39 : AX1B
      port map(A => \un1_state_12_2[4]\, B => 
        \un1_state_12_3_0[4]\, C => \addr_data_vector[2]\, Y => 
        N_40_i_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_24\ : OR2A
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => N_35_0);
    
    \state_ns_i_a2[1]\ : OR2A
      port map(A => update_and_sel_7(0), B => update_and_sel_7(1), 
        Y => N_83_i);
    
    un1_address_m23_m7_i_2 : NOR2B
      port map(A => \addr_data_vector[10]\, B => 
        \addr_data_vector[11]\, Y => m23_m7_i_2);
    
    \address_RNO[6]\ : MX2
      port map(A => \un1_address[6]\, B => addr_data_f0(6), S => 
        \state_0[0]_net_1\, Y => \address_7[6]\);
    
    \state_RNO[2]\ : AO1A
      port map(A => status_full_ack(0), B => N_84, C => N_80, Y
         => \state_ns[2]\);
    
    \address_RNIBG94[20]\ : MX2C
      port map(A => \addr_data_vector[20]\, B => 
        addr_data_vector_84, S => sel_data_1(1), Y => N_1313);
    
    \address_RNI7894[11]\ : MX2C
      port map(A => \addr_data_vector[11]\, B => 
        addr_data_vector_75, S => sel_data_1(1), Y => N_1318);
    
    \address_RNO[28]\ : MX2
      port map(A => \un1_address[28]\, B => addr_data_f0(28), S
         => \state[0]_net_1\, Y => \address_7[28]\);
    
    \address_RNO[11]\ : MX2
      port map(A => N_20_0_i_0, B => addr_data_f0(11), S => 
        \state_0[0]_net_1\, Y => \address_7[11]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_21\ : AO1C
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, C => N_30_0, Y => N_32);
    
    un1_address_m40_m6_0_a2_3 : NOR2B
      port map(A => \addr_data_vector[11]\, B => 
        \addr_data_vector[12]\, Y => m40_m6_0_a2_3);
    
    \FSM_SELECT_ADDRESS.state7_0_I_73\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => state7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_35\ : XNOR2
      port map(A => \un2_nb_send_next[5]\, B => 
        nb_burst_available(5), Y => \DWACT_BL_EQUAL_0_E[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_2\ : XNOR2
      port map(A => \un2_nb_send_next[6]\, B => 
        nb_burst_available(6), Y => \DWACT_BL_EQUAL_0_E_0[0]\);
    
    un1_address_m38 : AX1B
      port map(A => m23_m7_i, B => m37_m6_0_a2_4_i, C => 
        \addr_data_vector[23]\, Y => \un1_address[23]\);
    
    un1_address_m12 : AO13
      port map(A => N_5_0, B => address_0_sqmuxa, C => 
        \addr_data_vector[6]\, Y => N_13_0);
    
    un1_address_m59 : AX1
      port map(A => N_13_0, B => m40_m6_0_a2_7, C => 
        \addr_data_vector[24]\, Y => \un1_address[24]\);
    
    \update_r[0]\ : DFN1P0
      port map(D => update_and_sel_7(0), CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \update_r_i[0]\);
    
    un2_nb_send_next_I_5 : XOR2
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        Y => \un2_nb_send_next[1]\);
    
    \state_RNIBABE[1]\ : NOR2A
      port map(A => status_full_ack(0), B => N_85, Y => 
        \state_RNIBABE[1]_net_1\);
    
    un1_address_m40_m6_0_a2_6 : NOR3C
      port map(A => m40_m6_0_a2_3, B => m40_m6_0_a2_2, C => 
        m40_m6_0_a2_4, Y => m40_m6_0_a2_6);
    
    \address_RNO[17]\ : MX2
      port map(A => N_30_0_i_0, B => addr_data_f0(17), S => 
        \state[0]_net_1\, Y => \address_7[17]\);
    
    \address_RNO[5]\ : MX2
      port map(A => N_52_i_0, B => addr_data_f0(5), S => 
        \state_0[0]_net_1\, Y => \address_7[5]\);
    
    un1_address_m15 : OR3B
      port map(A => \addr_data_vector[7]\, B => 
        \addr_data_vector[8]\, C => N_13_0, Y => N_16_0);
    
    un1_address_m58 : AX1C
      port map(A => \addr_data_vector[21]\, B => N_36_0, C => 
        \addr_data_vector[22]\, Y => \un1_address[22]\);
    
    un2_nb_send_next_I_56 : XOR2
      port map(A => N_4, B => \nb_send[10]_net_1\, Y => 
        \un2_nb_send_next[10]\);
    
    un1_address_m26 : OR3B
      port map(A => \addr_data_vector[14]\, B => 
        \addr_data_vector[15]\, C => m23_m7_i, Y => N_27_0);
    
    un2_nb_send_next_I_41 : AND2
      port map(A => \nb_send[6]_net_1\, B => \nb_send[7]_net_1\, 
        Y => \DWACT_FINC_E[3]\);
    
    \address_RNO[3]\ : MX2
      port map(A => N_50_i_0, B => addr_data_f0(3), S => 
        \state_0[0]_net_1\, Y => \address_7[3]\);
    
    \address_RNO_4[31]\ : NOR2B
      port map(A => \addr_data_vector[28]\, B => 
        \addr_data_vector[29]\, Y => address_7_31_m6_e_2);
    
    \address[3]\ : DFN1C0
      port map(D => \address_7[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[3]\);
    
    un2_nb_send_next_I_34 : AND3
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        C => \nb_send[5]_net_1\, Y => \DWACT_FINC_E[2]\);
    
    un1_address_m64 : XOR2
      port map(A => N_46, B => \addr_data_vector[29]\, Y => 
        \un1_address[29]\);
    
    un1_address_m34 : XNOR2
      port map(A => N_34_0, B => \addr_data_vector[20]\, Y => 
        \un1_address[20]\);
    
    \address_RNO[30]\ : MX2
      port map(A => \un1_address[30]\, B => addr_data_f0(30), S
         => \state[0]_net_1\, Y => \address_7[30]\);
    
    \state_RNO_0[1]\ : OR2
      port map(A => status_full_ack(0), B => N_85, Y => 
        \state_ns_i_0[3]\);
    
    \nb_send[3]\ : DFN1E0C0
      port map(D => \nb_send_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[3]_net_1\);
    
    un1_address_m23_m7_i_1 : NOR2B
      port map(A => \addr_data_vector[8]\, B => 
        \addr_data_vector[9]\, Y => m23_m7_i_1);
    
    \address_RNIIVLA[0]\ : MX2C
      port map(A => \addr_data_vector[0]\, B => 
        addr_data_vector_64, S => sel_data_0(1), Y => N_1279);
    
    \FSM_SELECT_ADDRESS.state7_0_I_20\ : OR2A
      port map(A => nb_burst_available(10), B => 
        \un2_nb_send_next[10]\, Y => N_31);
    
    un1_address_m54 : AX1C
      port map(A => \addr_data_vector[12]\, B => N_21_0, C => 
        \addr_data_vector[13]\, Y => N_55_0_i_0);
    
    \address[7]\ : DFN1C0
      port map(D => \address_7[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[7]\);
    
    un2_nb_send_next_I_38 : XOR2
      port map(A => N_17, B => \nb_send[7]_net_1\, Y => 
        \un2_nb_send_next[7]\);
    
    \nb_send[5]\ : DFN1E0C0
      port map(D => \nb_send_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[5]_net_1\);
    
    un1_address_m3 : NOR3C
      port map(A => \addr_data_vector[3]\, B => N_2, C => 
        \addr_data_vector[4]\, Y => N_4_0);
    
    \nb_send_RNO[5]\ : NOR2B
      port map(A => \un2_nb_send_next[5]\, B => state7, Y => 
        \nb_send_5[5]\);
    
    \address_RNIDG94[21]\ : MX2C
      port map(A => \addr_data_vector[21]\, B => 
        addr_data_vector_85, S => sel_data_1(1), Y => N_1314);
    
    un1_address_m25 : AX1
      port map(A => m23_m7_i, B => \addr_data_vector[14]\, C => 
        \addr_data_vector[15]\, Y => N_26_0_i_0);
    
    \state[3]\ : DFN1C0
      port map(D => \state_RNO_1[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    
    \address_RNIFG94[22]\ : MX2C
      port map(A => \addr_data_vector[22]\, B => 
        addr_data_vector_86, S => sel_data_1(1), Y => N_1315);
    
    \update_r[1]\ : DFN1C0
      port map(D => update_and_sel_7(1), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \update_r[1]_net_1\);
    
    un1_address_m40_m6_0_a2_7 : NOR2A
      port map(A => m40_m6_0_a2_6, B => m37_m6_0_a2_4_i, Y => 
        m40_m6_0_a2_7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_17\ : OR2A
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, Y => N_28);
    
    \FSM_SELECT_ADDRESS.state7_0_I_43\ : AO1A
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => nb_burst_available(5), Y => 
        \ACT_LT2_E[2]\);
    
    \address_RNINHHB[4]\ : MX2C
      port map(A => \addr_data_vector[4]\, B => 
        addr_data_vector_68, S => sel_data(1), Y => N_1325);
    
    un1_address_m57 : XOR2
      port map(A => N_36_0, B => \addr_data_vector[21]\, Y => 
        \un1_address[21]\);
    
    un2_nb_send_next_I_8 : NOR2B
      port map(A => \nb_send[1]_net_1\, B => \nb_send[0]_net_1\, 
        Y => N_38);
    
    \address_RNING94[26]\ : MX2C
      port map(A => \addr_data_vector[26]\, B => 
        addr_data_vector_90, S => sel_data_1(1), Y => N_1305);
    
    \FSM_SELECT_ADDRESS.state7_0_I_23\ : AO1C
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), C => N_28, Y => N_34);
    
    \FSM_SELECT_ADDRESS.state7_0_I_26\ : OA1A
      port map(A => N_32, B => N_34, C => N_33, Y => N_37);
    
    \address_RNO[22]\ : MX2
      port map(A => \un1_address[22]\, B => addr_data_f0(22), S
         => \state[0]_net_1\, Y => \address_7[22]\);
    
    un2_nb_send_next_I_27 : AND2
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        Y => \DWACT_FINC_E[1]\);
    
    un1_address_m49 : XOR2
      port map(A => N_2, B => \addr_data_vector[3]\, Y => 
        N_50_i_0);
    
    \address[9]\ : DFN1C0
      port map(D => \address_7[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[9]\);
    
    \address_RNO[18]\ : MX2
      port map(A => \un1_address[18]\, B => addr_data_f0(18), S
         => \state[0]_net_1\, Y => \address_7[18]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \address_RNO[7]\ : MX2
      port map(A => N_1_i_0, B => addr_data_f0(7), S => 
        \state_0[0]_net_1\, Y => \address_7[7]\);
    
    un1_address_m23_m7_i_5 : NOR3C
      port map(A => m23_m7_i_2, B => m23_m7_i_1, C => m23_m7_i_3, 
        Y => m23_m7_i_5);
    
    \address[6]\ : DFN1C0
      port map(D => \address_7[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[6]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_59\ : OR2A
      port map(A => \un2_nb_send_next[3]\, B => 
        nb_burst_available(3), Y => \ACT_LT4_E[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_1\ : XNOR2
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => \DWACT_BL_EQUAL_0_E[4]\);
    
    \address_RNIRG94[28]\ : MX2C
      port map(A => \addr_data_vector[28]\, B => 
        addr_data_vector_92, S => sel_data_1(1), Y => N_1307);
    
    status_full_err_RNO : OR2
      port map(A => un1_state_5_i_0, B => N_84, Y => N_64);
    
    \state_0[0]\ : DFN1C0
      port map(D => \state_RNIBABE[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state_0[0]_net_1\);
    
    \address_RNO[8]\ : MX2
      port map(A => N_15_0_i_0, B => addr_data_f0(8), S => 
        \state_0[0]_net_1\, Y => \address_7[8]\);
    
    un2_nb_send_next_I_52 : XOR2
      port map(A => N_7, B => \nb_send[9]_net_1\, Y => 
        \un2_nb_send_next[9]\);
    
    \address[11]\ : DFN1C0
      port map(D => \address_7[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[11]\);
    
    \address[31]\ : DFN1C0
      port map(D => \address_7[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[31]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_55\ : OR2A
      port map(A => nb_burst_available(2), B => 
        \un2_nb_send_next[2]\, Y => \ACT_LT4_E[4]\);
    
    \state_RNIU3MB[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => un3_update_r, Y => 
        address_0_sqmuxa_0);
    
    un1_address_m56 : XNOR2
      port map(A => N_31_0, B => \addr_data_vector[18]\, Y => 
        \un1_address[18]\);
    
    \address_RNO[2]\ : MX2
      port map(A => N_40_i_0, B => addr_data_f0(2), S => 
        \state_0[0]_net_1\, Y => \address_7[2]\);
    
    \address_RNO[4]\ : MX2
      port map(A => N_51_i_0, B => addr_data_f0(4), S => 
        \state_0[0]_net_1\, Y => \address_7[4]\);
    
    un2_nb_send_next_I_19 : NOR2B
      port map(A => \nb_send[3]_net_1\, B => \DWACT_FINC_E[0]\, Y
         => N_30);
    
    \address_RNO[25]\ : MX2
      port map(A => \un1_address[25]\, B => addr_data_f0(25), S
         => \state[0]_net_1\, Y => \address_7[25]\);
    
    \address[21]\ : DFN1C0
      port map(D => \address_7[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[21]\);
    
    un1_address_m23_m7_i_3 : NOR3C
      port map(A => \addr_data_vector[7]\, B => 
        \addr_data_vector[13]\, C => \addr_data_vector[12]\, Y
         => m23_m7_i_3);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    un1_address_m62 : XOR2
      port map(A => N_44, B => \addr_data_vector[27]\, Y => 
        \un1_address[27]\);
    
    \address_RNIB894[13]\ : MX2C
      port map(A => \addr_data_vector[13]\, B => 
        addr_data_vector_77, S => sel_data_1(1), Y => N_1320);
    
    un1_address_m32 : AX1
      port map(A => N_31_0, B => \addr_data_vector[18]\, C => 
        \addr_data_vector[19]\, Y => \un1_address[19]\);
    
    un1_address_m12_e : OR2B
      port map(A => N_4_0, B => \addr_data_vector[5]\, Y => N_5_0);
    
    \address_RNO_5[31]\ : NOR2B
      port map(A => \addr_data_vector[26]\, B => 
        \addr_data_vector[27]\, Y => address_7_31_m6_e_1);
    
    un2_nb_send_next_I_9 : XOR2
      port map(A => N_38, B => \nb_send[2]_net_1\, Y => 
        \un2_nb_send_next[2]\);
    
    \state[1]\ : DFN1C0
      port map(D => \state_RNO_0[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state[1]_net_1\);
    
    \address[17]\ : DFN1C0
      port map(D => \address_7[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[17]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_52\ : OR2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[1]\);
    
    un1_address_m65 : AX1C
      port map(A => \addr_data_vector[29]\, B => N_46, C => 
        \addr_data_vector[30]\, Y => \un1_address[30]\);
    
    un1_address_m35 : NOR2A
      port map(A => \addr_data_vector[20]\, B => N_34_0, Y => 
        N_36_0);
    
    un1_address_m52 : XNOR2
      port map(A => N_13_0, B => \addr_data_vector[7]\, Y => 
        N_1_i_0);
    
    \address_RNINFMA[2]\ : MX2C
      port map(A => \addr_data_vector[2]\, B => 
        addr_data_vector_66, S => sel_data_1(1), Y => N_1323);
    
    \address[27]\ : DFN1C0
      port map(D => \address_7[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[27]\);
    
    \state_RNO[3]\ : NOR2B
      port map(A => \state[4]_net_1\, B => N_83_i, Y => 
        \state_RNO_1[3]\);
    
    un1_address_m21 : XOR2
      port map(A => N_21_0, B => \addr_data_vector[12]\, Y => 
        N_22_0_i_0);
    
    \nb_send_RNO[4]\ : NOR2B
      port map(A => \un2_nb_send_next[4]\, B => state7, Y => 
        \nb_send_5[4]\);
    
    \nb_send_RNO[10]\ : NOR2B
      port map(A => \un2_nb_send_next[10]\, B => state7, Y => 
        \nb_send_5[10]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_18\ : OR2A
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => N_29);
    
    \address_RNIGO94[30]\ : MX2C
      port map(A => \addr_data_vector[30]\, B => 
        addr_data_vector_94, S => sel_data_0(1), Y => N_1295);
    
    un1_address_m55 : XNOR2
      port map(A => m23_m7_i, B => \addr_data_vector[14]\, Y => 
        N_56_0_i_0);
    
    \address_RNO[31]\ : MX2C
      port map(A => \address_RNO_0_0[31]\, B => 
        \address_RNO_1_0[31]\, S => \address_RNO_2_0[31]\, Y => 
        \address_7[31]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_61\ : AOI1A
      port map(A => \ACT_LT4_E[3]\, B => \ACT_LT4_E[6]\, C => 
        \ACT_LT4_E[10]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_34\ : XNOR2
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), Y => \DWACT_BL_EQUAL_0_E[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_6\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E_0[0]\, B => 
        \DWACT_BL_EQUAL_0_E_0[1]\, C => \DWACT_BL_EQUAL_0_E[2]\, 
        Y => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\);
    
    \address_RNO[12]\ : MX2
      port map(A => N_22_0_i_0, B => addr_data_f0(12), S => 
        \state_0[0]_net_1\, Y => \address_7[12]\);
    
    \update_r_RNIVJV4_0[0]\ : OR2
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => \un1_state_12_3_0[4]\);
    
    un2_nb_send_next_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \nb_send[6]_net_1\, Y => N_17);
    
    un2_nb_send_next_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_12);
    
    \FSM_SELECT_ADDRESS.state7_0_I_3\ : XNOR2
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => \DWACT_BL_EQUAL_0_E[2]\);
    
    status_full_RNO : OR2
      port map(A => \state[2]_net_1\, B => N_80, Y => 
        un1_state_11);
    
    \address_RNIJG94[24]\ : MX2C
      port map(A => \addr_data_vector[24]\, B => 
        addr_data_vector_88, S => sel_data_1(1), Y => N_1303);
    
    \address[1]\ : DFN1E1C0
      port map(D => addr_data_f0(1), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        \addr_data_vector[1]\);
    
    \status_full\ : DFN1E1C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_11, Q => status_full(0));
    
    un1_address_m63 : AX1C
      port map(A => \addr_data_vector[27]\, B => N_44, C => 
        \addr_data_vector[28]\, Y => \un1_address[28]\);
    
    un1_address_m33 : OR3B
      port map(A => \addr_data_vector[18]\, B => 
        \addr_data_vector[19]\, C => N_31_0, Y => N_34_0);
    
    \state_RNIA6SP8_0[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => state7, Y => N_80);
    
    un2_nb_send_next_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    \address_RNO[20]\ : MX2
      port map(A => \un1_address[20]\, B => addr_data_f0(20), S
         => \state[0]_net_1\, Y => \address_7[20]\);
    
    \nb_send[8]\ : DFN1E0C0
      port map(D => \nb_send_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[8]_net_1\);
    
    \address_RNIL894[18]\ : MX2C
      port map(A => \addr_data_vector[18]\, B => 
        addr_data_vector_82, S => sel_data_1(1), Y => N_1311);
    
    un1_address_m53 : AX1
      port map(A => N_16_0, B => \addr_data_vector[9]\, C => 
        \addr_data_vector[10]\, Y => N_54_0_i_0);
    
    un1_address_m40_m6_0_a2_1 : NOR2B
      port map(A => \addr_data_vector[7]\, B => 
        \addr_data_vector[8]\, Y => m40_m6_0_a2_1);
    
    \address_RNO_3[31]\ : NOR3C
      port map(A => \addr_data_vector[25]\, B => 
        \addr_data_vector[30]\, C => address_7_31_m6_e_1, Y => 
        address_7_31_m6_e_3);
    
    un1_address_m37_m6_0_a2_4_4 : NOR3C
      port map(A => \addr_data_vector[14]\, B => 
        \addr_data_vector[22]\, C => \addr_data_vector[21]\, Y
         => m37_m6_0_a2_4_4);
    
    \nb_send[1]\ : DFN1E0C0
      port map(D => \nb_send_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_60\ : AOI1A
      port map(A => \ACT_LT4_E[7]\, B => \ACT_LT4_E[8]\, C => 
        \ACT_LT4_E[5]\, Y => \ACT_LT4_E[10]\);
    
    \state_RNO_1[4]\ : OR3A
      port map(A => \state_0[0]_net_1\, B => \state[3]_net_1\, C
         => \state[2]_net_1\, Y => N_78);
    
    \address_RNO[15]\ : MX2
      port map(A => N_26_0_i_0, B => addr_data_f0(15), S => 
        \state_0[0]_net_1\, Y => \address_7[15]\);
    
    un2_nb_send_next_I_20 : XOR2
      port map(A => N_30, B => \nb_send[4]_net_1\, Y => 
        \un2_nb_send_next[4]\);
    
    un1_address_m37_m6_0_a2_4_5 : NOR3C
      port map(A => \addr_data_vector[16]\, B => 
        \addr_data_vector[15]\, C => m37_m6_0_a2_4_2, Y => 
        m37_m6_0_a2_4_5);
    
    \FSM_SELECT_ADDRESS.state7_0_I_68\ : AO1
      port map(A => \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, B => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, C => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, Y => 
        \DWACT_COMP0_E[2]\);
    
    un2_nb_send_next_I_16 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_dma_send_16word is

    port( un7_dmain        : out   std_logic_vector(66 to 66);
          data_address     : in    std_logic_vector(31 downto 0);
          Store            : out   std_logic;
          Fault            : in    std_logic;
          un1_data_send_ok : out   std_logic;
          Request_0        : in    std_logic;
          N_1011           : out   std_logic;
          Lock_0           : in    std_logic;
          N_1013           : out   std_logic;
          N_957            : out   std_logic;
          N_956            : out   std_logic;
          N_955            : out   std_logic;
          N_954            : out   std_logic;
          N_953            : out   std_logic;
          N_952            : out   std_logic;
          N_951            : out   std_logic;
          N_964            : out   std_logic;
          N_963            : out   std_logic;
          N_962            : out   std_logic;
          N_961            : out   std_logic;
          N_960            : out   std_logic;
          time_select      : in    std_logic;
          N_959            : out   std_logic;
          N_958            : out   std_logic;
          N_971            : out   std_logic;
          N_970            : out   std_logic;
          N_969            : out   std_logic;
          N_968            : out   std_logic;
          N_967            : out   std_logic;
          N_966            : out   std_logic;
          N_965            : out   std_logic;
          N_978            : out   std_logic;
          N_977            : out   std_logic;
          N_976            : out   std_logic;
          N_975            : out   std_logic;
          N_974            : out   std_logic;
          N_973            : out   std_logic;
          N_972            : out   std_logic;
          N_950            : out   std_logic;
          N_949            : out   std_logic;
          N_948            : out   std_logic;
          time_select_0    : in    std_logic;
          N_947            : out   std_logic;
          N_249            : out   std_logic;
          Grant            : in    std_logic;
          Ready            : in    std_logic;
          data_send        : in    std_logic;
          OKAY             : in    std_logic;
          N_200            : out   std_logic;
          HRESETn_c        : in    std_logic;
          HCLK_c           : in    std_logic
        );

end lpp_dma_send_16word;

architecture DEF_ARCH of lpp_dma_send_16word is 

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \state_0[5]_net_1\, N_4, N_198_0, N_509, N_344, 
        N_154_0, N_241, N_235, N_242, N_202_0, m74_0, 
        \data_counter[30]_net_1\, \data_counter[29]_net_1\, 
        ADD_32x32_fast_I129_un1_Y_14, ADD_32x32_fast_I129_un1_Y_9, 
        ADD_32x32_fast_I129_un1_Y_8, ADD_32x32_fast_I129_un1_Y_13, 
        ADD_32x32_fast_I129_un1_Y_5, ADD_32x32_fast_I129_un1_Y_4, 
        ADD_32x32_fast_I129_un1_Y_11, \grant_counter[27]_net_1\, 
        \grant_counter[26]_net_1\, ADD_32x32_fast_I129_un1_Y_7, 
        \grant_counter[19]_net_1\, \grant_counter[18]_net_1\, 
        ADD_32x32_fast_I129_un1_Y_3, \grant_counter[15]_net_1\, 
        \grant_counter[14]_net_1\, ADD_32x32_fast_I129_un1_Y_1, 
        \grant_counter[28]_net_1\, \grant_counter[29]_net_1\, 
        \grant_counter[24]_net_1\, \grant_counter[25]_net_1\, 
        \grant_counter[22]_net_1\, \grant_counter[23]_net_1\, 
        \grant_counter[20]_net_1\, \grant_counter[21]_net_1\, 
        \grant_counter[16]_net_1\, \grant_counter[17]_net_1\, 
        m43_m6_0_a2_6, \grant_counter[13]_net_1\, 
        \grant_counter[12]_net_1\, m43_m6_0_a2_4, m43_m6_0_a2_5, 
        \grant_counter[9]_net_1\, \grant_counter[8]_net_1\, 
        m43_m6_0_a2_2, \grant_counter[7]_net_1\, 
        \grant_counter[6]_net_1\, \grant_counter[10]_net_1\, 
        \grant_counter[11]_net_1\, \data_counter_8_i_0[0]\, N_508, 
        N_338_1, N_337, \grant_counter_0_i_0[4]\, N_246, 
        un1_hresetn_inv_i_0, ADD_32x32_fast_I129_un1_Y_14_0, 
        ADD_32x32_fast_I129_un1_Y_9_0, 
        ADD_32x32_fast_I129_un1_Y_8_0, 
        ADD_32x32_fast_I129_un1_Y_13_0, 
        ADD_32x32_fast_I129_un1_Y_5_0, 
        ADD_32x32_fast_I129_un1_Y_4_0, 
        ADD_32x32_fast_I129_un1_Y_11_0, \data_counter[27]_net_1\, 
        \data_counter[26]_net_1\, ADD_32x32_fast_I129_un1_Y_7_0, 
        \data_counter[19]_net_1\, \data_counter[18]_net_1\, 
        ADD_32x32_fast_I129_un1_Y_3_0, \data_counter[15]_net_1\, 
        \data_counter[14]_net_1\, ADD_32x32_fast_I129_un1_Y_1_0, 
        \data_counter[28]_net_1\, \data_counter[24]_net_1\, 
        \data_counter[25]_net_1\, \data_counter[22]_net_1\, 
        \data_counter[23]_net_1\, \data_counter[20]_net_1\, 
        \data_counter[21]_net_1\, \data_counter[16]_net_1\, 
        \data_counter[17]_net_1\, m28_m6_5, \state[3]_net_1\, 
        m28_m6_4, m28_m6_1, m28_m6_0, m28_m6_2, 
        \data_counter[0]_net_1\, \state[0]_net_1\, 
        \data_counter[2]_net_1\, \data_counter[3]_net_1\, 
        \data_counter[13]_net_1\, \data_counter[1]_net_1\, 
        \grant_counter_0_0_0[0]\, \grant_counter[0]_net_1\, 
        un1_state_2_i_o2_0, \state[1]_net_1\, \state[2]_net_1\, 
        \state_ns_i_a2_i_0_0[0]\, un1_state_7_i_a4_0_1, N_518_1, 
        un1_state_5_i_o2_30, un1_state_5_i_o2_25, 
        un1_state_5_i_o2_24, un1_state_5_i_o2_29, 
        un1_state_5_i_o2_21, un1_state_5_i_o2_20, 
        un1_state_5_i_o2_27, un1_state_5_i_o2_13, 
        un1_state_5_i_o2_12, un1_state_5_i_o2_23, 
        un1_state_5_i_o2_5, un1_state_5_i_o2_4, 
        un1_state_5_i_o2_19, un1_state_5_i_o2_1, 
        un1_state_5_i_o2_0, un1_state_5_i_o2_17, 
        un1_state_5_i_o2_15, un1_state_5_i_o2_11, 
        un1_state_5_i_o2_9, un1_state_5_i_o2_7, 
        un1_state_5_i_o2_3, \data_counter[5]_net_1\, 
        \data_counter[4]_net_1\, \data_counter[10]_net_1\, 
        \data_counter[11]_net_1\, \data_counter[8]_net_1\, 
        \data_counter[9]_net_1\, \data_counter[6]_net_1\, 
        \data_counter[7]_net_1\, \data_counter[31]_net_1\, 
        \data_counter[12]_net_1\, \state_ns_i_a2_0_i_o2_29[3]\, 
        \state_ns_i_a2_0_i_o2_21[3]\, 
        \state_ns_i_a2_0_i_o2_20[3]\, 
        \state_ns_i_a2_0_i_o2_27[3]\, 
        \state_ns_i_a2_0_i_o2_22[3]\, 
        \state_ns_i_a2_0_i_o2_23[3]\, 
        \state_ns_i_a2_0_i_o2_25[3]\, \state_ns_i_a2_0_i_o2_5[3]\, 
        \state_ns_i_a2_0_i_o2_4[3]\, \state_ns_i_a2_0_i_o2_19[3]\, 
        \state_ns_i_a2_0_i_o2_24[3]\, \state_ns_i_a2_0_i_o2_3[3]\, 
        \state_ns_i_a2_0_i_o2_2[3]\, \state_ns_i_a2_0_i_o2_16[3]\, 
        \state_ns_i_a2_0_i_o2_15[3]\, 
        \state_ns_i_a2_0_i_o2_13[3]\, 
        \state_ns_i_a2_0_i_o2_11[3]\, \state_ns_i_a2_0_i_o2_9[3]\, 
        \state_ns_i_a2_0_i_o2_6[3]\, \state_ns_i_a2_0_i_o2_7[3]\, 
        \state_ns_i_a2_0_i_o2_1[3]\, \grant_counter[4]_net_1\, 
        \grant_counter[31]_net_1\, \grant_counter[2]_net_1\, 
        \grant_counter[3]_net_1\, \grant_counter[1]_net_1\, 
        \grant_counter[5]_net_1\, \grant_counter[30]_net_1\, 
        m27_m6_0_a2_4_5, m27_m6_0_a2_4_2, m27_m6_0_a2_4_4, 
        m27_m6_0_a2_4_3, N_75, N_72, I129_un1_Y, N623, 
        \grant_counter_RNO[0]_net_1\, N_89, N_19_0, N_346, N_243, 
        \state[4]_net_1\, N_194_i_0, N_522, Burst, N_526, N_339, 
        N_186, N_336, \un1_state_4_i_i[31]\, N_75_0, N_72_0, 
        m27_m6_0_a2_4, N_44, N_21_0, N623_0, N_28_0, N_19_0_0, 
        N_22_0, N_23_0, N_24_0, N_25_0, N_26_0, N_27_0, N_28_0_0, 
        \un1_hresetn_inv_2_i[26]\, \un1_hresetn_inv_2_i[15]\, 
        N_48, \un1_hresetn_inv_2_i[13]\, N_52, 
        \un1_hresetn_inv_2_i[11]\, N_56, \un1_hresetn_inv_2_i[9]\, 
        N_60, \un1_hresetn_inv_2_i[7]\, N_64, 
        \un1_hresetn_inv_2_i[5]\, N_68, \un1_hresetn_inv_2_i[3]\, 
        N_23_0_0, N_22_0_0, N_24_0_0, N_25_0_0, N_26_0_0, 
        N_27_0_0, N_45, N_46, N_48_0, N_50, N_52_0, N_54, N_56_0, 
        N_58, N_60_0, N_62, N_64_0, N_66, N_68_0, 
        \un1_state_4_i[17]\, \data_counter_8[7]\, 
        \data_counter_8[8]\, \data_counter_8[9]\, 
        \data_counter_8[10]\, \data_counter_8[11]\, 
        \data_counter_8[12]\, \data_counter_8[13]\, 
        \data_counter_8[14]\, \data_counter_8[15]\, 
        \data_counter_8[16]\, \data_counter_8[17]\, 
        \data_counter_8[18]\, \data_counter_8[19]\, 
        \data_counter_8[20]\, \data_counter_8[21]\, N_198, 
        \data_counter_8[22]\, \data_counter_8[23]\, 
        \data_counter_8[24]\, \data_counter_8[25]\, 
        \data_counter_8[26]\, N_13, N_15, N_17, N_19, N_21, N_23, 
        N_25, N_27, N_29, N_31, N_33, N_35, N_43, N_45_0, N_47, 
        N_49, N_51, N_53, N_55, \state[5]_net_1\, N_57, N_59, 
        N_61, N_63, N_65, N_67, N_69, N_71, N_73, N_75_1, N_77, 
        N_79, N_81, N_91, N_93, N_95, N_97, N_99, N_101, N_103, 
        N_105, N_107, N_109, N_111, N_113, N_115, N_117, N_119, 
        N_202, N_121, N_123, N_125, N_127, N_129, N_131, N_133, 
        N_135, N_137, N_139, N_141, N_143, \N_200\, \Address[0]\, 
        \Address[1]\, \Address[2]\, \Address[3]\, \Address[25]\, 
        \Address[26]\, \Address[27]\, \Address[28]\, 
        \Address[29]\, \Address[30]\, \Address[31]\, 
        \Address[18]\, \Address[19]\, \Address[20]\, 
        \Address[21]\, \Address[22]\, \Address[23]\, 
        \Address[24]\, \Address[11]\, \Address[12]\, 
        \Address[13]\, \Address[14]\, \Address[15]\, 
        \Address[16]\, \Address[17]\, \Address[4]\, \Address[5]\, 
        \Address[6]\, \Address[7]\, \Address[8]\, \Address[9]\, 
        \Address[10]\, Lock, Request, N_84, Request_5, N_32_0_i_0, 
        N_17_0, \grant_counter_RNO[2]_net_1\, N_513, N_146, N_516, 
        N_151, data_send_ok, data_send_ko, 
        \grant_counter_RNO[3]_net_1\, N_33_0_i_0, 
        \grant_counter_RNO[1]_net_1\, N_31_0_i_0, 
        \state_RNO_0[0]_net_1\, \state_RNO[0]_net_1\, 
        \state_RNO[3]_net_1\, N_154, N_192, \un1_state_4_i[28]\, 
        N_190, \un1_state_4_i[29]\, N_188, \un1_state_4_i[30]\, 
        N_156, N_348, \data_counter_8[31]\, \data_counter_8[30]\, 
        \un1_state_4_i[1]\, \data_counter_8[29]\, 
        \data_counter_8[28]\, N_70, \data_counter_8[27]\, 
        \data_counter_8[6]\, N_21_0_0, \data_counter_8[5]\, 
        N_20_0, \data_counter_8[4]\, N_510, N_18_0, N_16_0, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    N_200 <= \N_200\;

    un1_hresetn_inv_2_m66 : AX1E
      port map(A => \grant_counter[25]_net_1\, B => N_64, C => 
        \grant_counter[26]_net_1\, Y => \un1_hresetn_inv_2_i[5]\);
    
    \state_RNIK8SG_1[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => OKAY, Y => N_249);
    
    \DMAIn.Address[7]\ : DFN1E1C0
      port map(D => N_27, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[7]\);
    
    \state[0]\ : DFN1C0
      port map(D => \state_RNO[0]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[0]_net_1\);
    
    un1_state_4_m28_m6_4 : NOR3C
      port map(A => m28_m6_1, B => m28_m6_0, C => m28_m6_2, Y => 
        m28_m6_4);
    
    \data_counter_RNIMF78[4]\ : NOR3A
      port map(A => un1_state_5_i_o2_3, B => 
        \data_counter[5]_net_1\, C => \data_counter[4]_net_1\, Y
         => un1_state_5_i_o2_17);
    
    \data_counter_RNO[31]\ : XA1C
      port map(A => \data_counter[31]_net_1\, B => N_75_0, C => 
        N_198, Y => \data_counter_8[31]\);
    
    un1_state_4_m51 : NOR2B
      port map(A => N_50, B => \data_counter[18]_net_1\, Y => 
        N_52_0);
    
    \data_counter_RNO[2]\ : AOI1B
      port map(A => \un1_state_4_i[29]\, B => N_344, C => N_509, 
        Y => N_190);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_3 : NOR2B
      port map(A => \grant_counter[20]_net_1\, B => 
        \grant_counter[21]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_3);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y : NOR2B
      port map(A => ADD_32x32_fast_I129_un1_Y_14, B => N623, Y
         => I129_un1_Y);
    
    \data_counter_RNO[18]\ : XA1B
      port map(A => \data_counter[18]_net_1\, B => N_50, C => 
        N_198_0, Y => \data_counter_8[18]\);
    
    un1_state_4_m17 : NOR3C
      port map(A => \data_counter[1]_net_1\, B => N_16_0, C => 
        \data_counter[2]_net_1\, Y => N_18_0);
    
    \grant_counter_RNO[5]\ : NOR2A
      port map(A => N_202_0, B => \un1_hresetn_inv_2_i[26]\, Y
         => N_91);
    
    un1_state_4_m49 : NOR2B
      port map(A => N_48_0, B => \data_counter[17]_net_1\, Y => 
        N_50);
    
    un1_state_4_m28_m6_2 : NOR2A
      port map(A => \data_counter[0]_net_1\, B => 
        \state[0]_net_1\, Y => m28_m6_2);
    
    \DMAIn.Address_RNIJIRJ[25]\ : MX2
      port map(A => \Address[25]\, B => data_address(25), S => 
        time_select_0, Y => N_972);
    
    \DMAIn.Address_RNI54FJ[14]\ : MX2
      port map(A => \Address[14]\, B => data_address(14), S => 
        time_select, Y => N_961);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_5 : NOR2B
      port map(A => \data_counter[24]_net_1\, B => 
        \data_counter[25]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_5_0);
    
    \grant_counter_RNO[26]\ : NOR2A
      port map(A => N_202, B => \un1_hresetn_inv_2_i[5]\, Y => 
        N_133);
    
    \DMAIn.Address_RNO[20]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(20), Y
         => N_59);
    
    \DMAIn.Address_RNIEF261[5]\ : MX2
      port map(A => \Address[5]\, B => data_address(5), S => 
        time_select, Y => N_952);
    
    \grant_counter[0]\ : DFN1
      port map(D => \grant_counter_RNO[0]_net_1\, CLK => HCLK_c, 
        Q => \grant_counter[0]_net_1\);
    
    \DMAIn.Address[6]\ : DFN1E1C0
      port map(D => N_25, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[6]\);
    
    \DMAIn.Address_RNI3IKI[13]\ : MX2
      port map(A => \Address[13]\, B => data_address(13), S => 
        time_select, Y => N_960);
    
    \DMAIn.Address_RNIL0M41[0]\ : MX2
      port map(A => \Address[0]\, B => data_address(0), S => 
        time_select_0, Y => N_947);
    
    un1_state_4_m53 : NOR2B
      port map(A => N_52_0, B => \data_counter[19]_net_1\, Y => 
        N_54);
    
    \grant_counter[20]\ : DFN1
      port map(D => N_121, CLK => HCLK_c, Q => 
        \grant_counter[20]_net_1\);
    
    \DMAIn.Address_RNO[27]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(27), Y
         => N_73);
    
    un1_state_4_m27_m6_0_a2_4_4 : NOR3C
      port map(A => \data_counter[4]_net_1\, B => 
        \data_counter[12]_net_1\, C => \data_counter[11]_net_1\, 
        Y => m27_m6_0_a2_4_4);
    
    \data_counter_RNO[14]\ : NOR2
      port map(A => \un1_state_4_i[17]\, B => N_198_0, Y => 
        \data_counter_8[14]\);
    
    \data_counter_RNO[21]\ : XA1B
      port map(A => \data_counter[21]_net_1\, B => N_56_0, C => 
        N_198, Y => \data_counter_8[21]\);
    
    \data_counter_RNIN6PF[31]\ : NOR2
      port map(A => \data_counter[31]_net_1\, B => 
        \data_counter[12]_net_1\, Y => un1_state_5_i_o2_0);
    
    \DMAIn.Address[2]\ : DFN1E1C0
      port map(D => N_17, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[2]\);
    
    \DMAIn.Address[28]\ : DFN1E1C0
      port map(D => N_75_1, CLK => HCLK_c, CLR => HRESETn_c, E
         => N_154, Q => \Address[28]\);
    
    un1_state_4_m19 : NOR2B
      port map(A => N_19_0_0, B => \data_counter[4]_net_1\, Y => 
        N_20_0);
    
    \grant_counter[26]\ : DFN1
      port map(D => N_133, CLK => HCLK_c, Q => 
        \grant_counter[26]_net_1\);
    
    \grant_counter[29]\ : DFN1
      port map(D => N_139, CLK => HCLK_c, Q => 
        \grant_counter[29]_net_1\);
    
    \grant_counter[1]\ : DFN1
      port map(D => \grant_counter_RNO[1]_net_1\, CLK => HCLK_c, 
        Q => \grant_counter[1]_net_1\);
    
    \data_counter[16]\ : DFN1C0
      port map(D => \data_counter_8[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[16]_net_1\);
    
    \data_counter[13]\ : DFN1C0
      port map(D => \data_counter_8[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[13]_net_1\);
    
    un1_state_4_m74 : OR2B
      port map(A => m74_0, B => N_72_0, Y => N_75_0);
    
    un1_hresetn_inv_2_m21 : NOR2B
      port map(A => N_21_0, B => \grant_counter[6]_net_1\, Y => 
        N_22_0);
    
    \state_0[5]\ : DFN1P0
      port map(D => N_4, CLK => HCLK_c, PRE => HRESETn_c, Q => 
        \state_0[5]_net_1\);
    
    \DMAIn.Address[29]\ : DFN1E1C0
      port map(D => N_77, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[29]\);
    
    \state_RNIV6P14[3]\ : OR2A
      port map(A => N_526, B => N_242, Y => N_156);
    
    \grant_counter_RNO[3]\ : AO1
      port map(A => N_33_0_i_0, B => N_202, C => N_513, Y => 
        \grant_counter_RNO[3]_net_1\);
    
    \grant_counter_RNIP43F[6]\ : NOR2
      port map(A => \grant_counter[6]_net_1\, B => 
        \grant_counter[7]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_4[3]\);
    
    un1_hresetn_inv_2_m20 : NOR3C
      port map(A => \grant_counter[4]_net_1\, B => N_19_0, C => 
        \grant_counter[5]_net_1\, Y => N_21_0);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_9 : NOR3C
      port map(A => \data_counter[19]_net_1\, B => 
        \data_counter[18]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_3_0, Y => 
        ADD_32x32_fast_I129_un1_Y_9_0);
    
    \grant_counter_RNIC1Q[18]\ : NOR3A
      port map(A => \state_ns_i_a2_0_i_o2_11[3]\, B => 
        \grant_counter[19]_net_1\, C => \grant_counter[18]_net_1\, 
        Y => \state_ns_i_a2_0_i_o2_21[3]\);
    
    \grant_counter_RNIBSC[10]\ : NOR2
      port map(A => \grant_counter[10]_net_1\, B => 
        \grant_counter[11]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_6[3]\);
    
    \grant_counter_RNO[16]\ : NOR2A
      port map(A => N_202_0, B => \un1_hresetn_inv_2_i[15]\, Y
         => N_113);
    
    un1_hresetn_inv_2_m23 : NOR2B
      port map(A => N_23_0, B => \grant_counter[8]_net_1\, Y => 
        N_24_0);
    
    \data_counter[11]\ : DFN1C0
      port map(D => \data_counter_8[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[11]_net_1\);
    
    \data_counter_RNIMDJV[22]\ : NOR3A
      port map(A => un1_state_5_i_o2_11, B => 
        \data_counter[23]_net_1\, C => \data_counter[22]_net_1\, 
        Y => un1_state_5_i_o2_21);
    
    \data_counter_RNI4TP71[4]\ : NOR3C
      port map(A => un1_state_5_i_o2_1, B => un1_state_5_i_o2_0, 
        C => un1_state_5_i_o2_17, Y => un1_state_5_i_o2_24);
    
    \data_counter[8]\ : DFN1C0
      port map(D => \data_counter_8[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[8]_net_1\);
    
    \grant_counter_RNO[4]\ : XA1B
      port map(A => \grant_counter[4]_net_1\, B => N_19_0, C => 
        \grant_counter_0_i_0[4]\, Y => N_89);
    
    \DMAIn.Address[1]\ : DFN1E1C0
      port map(D => N_15, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[1]\);
    
    \DMAIn.Address[13]\ : DFN1E1C0
      port map(D => N_45_0, CLK => HCLK_c, CLR => HRESETn_c, E
         => N_154_0, Q => \Address[13]\);
    
    \state_RNIRGVK7[0]\ : OR2A
      port map(A => N_348, B => N_235, Y => N_344);
    
    \state_RNI97HH[3]\ : MX2B
      port map(A => \state[5]_net_1\, B => Fault, S => 
        \state[3]_net_1\, Y => N_242);
    
    \grant_counter_RNIH42F[3]\ : NOR2B
      port map(A => \grant_counter[2]_net_1\, B => 
        \grant_counter[3]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_3[3]\);
    
    \DMAIn.Address[30]\ : DFN1E1C0
      port map(D => N_79, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[30]\);
    
    \DMAIn.Address_RNO[0]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(0), Y
         => N_13);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_8 : NOR3C
      port map(A => \grant_counter[15]_net_1\, B => 
        \grant_counter[14]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_1, Y => 
        ADD_32x32_fast_I129_un1_Y_8);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_5 : NOR2B
      port map(A => \grant_counter[24]_net_1\, B => 
        \grant_counter[25]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_5);
    
    un1_hresetn_inv_2_m26 : NOR2B
      port map(A => N_26_0, B => \grant_counter[11]_net_1\, Y => 
        N_27_0);
    
    \DMAIn.Address_RNO[10]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(10), Y
         => N_33);
    
    \DMAIn.Address_RNO[5]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(5), Y
         => N_23);
    
    send_ok : DFN1E1C0
      port map(D => \state[0]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_146, Q => data_send_ok);
    
    \grant_counter_RNO[9]\ : XA1
      port map(A => \grant_counter[9]_net_1\, B => N_24_0, C => 
        N_202_0, Y => N_99);
    
    \data_counter_RNI5VQF[28]\ : NOR2
      port map(A => \data_counter[28]_net_1\, B => 
        \data_counter[29]_net_1\, Y => un1_state_5_i_o2_13);
    
    \DMAIn.Address[31]\ : DFN1E1C0
      port map(D => N_81, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[31]\);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_11 : NOR3C
      port map(A => \grant_counter[27]_net_1\, B => 
        \grant_counter[26]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_7, Y => 
        ADD_32x32_fast_I129_un1_Y_11);
    
    \grant_counter_RNIC1GF[31]\ : NOR3A
      port map(A => \state_ns_i_a2_0_i_o2_1[3]\, B => 
        \grant_counter[4]_net_1\, C => \grant_counter[31]_net_1\, 
        Y => \state_ns_i_a2_0_i_o2_16[3]\);
    
    \DMAIn.Address_RNIMP5I[11]\ : MX2
      port map(A => \Address[11]\, B => data_address(11), S => 
        time_select_0, Y => N_958);
    
    \grant_counter[25]\ : DFN1
      port map(D => N_131, CLK => HCLK_c, Q => 
        \grant_counter[25]_net_1\);
    
    \DMAIn.Address_RNO[17]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(17), Y
         => N_53);
    
    un1_state_4_m18 : NOR2B
      port map(A => N_18_0, B => \data_counter[3]_net_1\, Y => 
        N_19_0_0);
    
    un1_state_4_m55 : NOR2B
      port map(A => N_54, B => \data_counter[20]_net_1\, Y => 
        N_56_0);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_1 : NOR2B
      port map(A => \data_counter[16]_net_1\, B => 
        \data_counter[17]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_1_0);
    
    un1_hresetn_inv_2_m71 : NOR3C
      port map(A => \grant_counter[27]_net_1\, B => N_68, C => 
        \grant_counter[28]_net_1\, Y => N_72);
    
    \state[4]\ : DFN1C0
      port map(D => N_84, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[4]_net_1\);
    
    \grant_counter_RNO[6]\ : XA1
      port map(A => \grant_counter[6]_net_1\, B => N_21_0, C => 
        N_202_0, Y => N_93);
    
    \data_counter_RNO[22]\ : XA1B
      port map(A => \data_counter[22]_net_1\, B => N_58, C => 
        N_198, Y => \data_counter_8[22]\);
    
    un1_hresetn_inv_2_m70 : AX1E
      port map(A => \grant_counter[27]_net_1\, B => N_68, C => 
        \grant_counter[28]_net_1\, Y => \un1_hresetn_inv_2_i[3]\);
    
    \DMAIn.Address_RNO[28]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(28), Y
         => N_75_1);
    
    \DMAIn.Address_RNI09N41[2]\ : MX2
      port map(A => \Address[2]\, B => data_address(2), S => 
        time_select_0, Y => N_949);
    
    \data_counter_RNITN34[6]\ : NOR2
      port map(A => \data_counter[6]_net_1\, B => 
        \data_counter[7]_net_1\, Y => un1_state_5_i_o2_3);
    
    \DMAIn.Address_RNIUHKI[12]\ : MX2
      port map(A => \Address[12]\, B => data_address(12), S => 
        time_select, Y => N_959);
    
    \data_counter_RNI1FQF[26]\ : NOR2
      port map(A => \data_counter[26]_net_1\, B => 
        \data_counter[27]_net_1\, Y => un1_state_5_i_o2_12);
    
    \grant_counter_RNO[20]\ : NOR2A
      port map(A => N_202, B => \un1_hresetn_inv_2_i[11]\, Y => 
        N_121);
    
    un1_state_4_m21 : NOR2B
      port map(A => N_21_0_0, B => \data_counter[6]_net_1\, Y => 
        N_22_0_0);
    
    \grant_counter_RNITK3F[8]\ : NOR2
      port map(A => \grant_counter[8]_net_1\, B => 
        \grant_counter[9]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_5[3]\);
    
    un1_hresetn_inv_2_m59 : NOR3C
      port map(A => \grant_counter[21]_net_1\, B => N_56, C => 
        \grant_counter[22]_net_1\, Y => N_60);
    
    \data_counter_RNIJJIB3[4]\ : NOR3B
      port map(A => un1_state_5_i_o2_25, B => un1_state_5_i_o2_24, 
        C => OKAY, Y => un1_state_5_i_o2_30);
    
    \grant_counter_RNO[22]\ : NOR2A
      port map(A => N_202, B => \un1_hresetn_inv_2_i[9]\, Y => 
        N_125);
    
    un1_state_4_m22 : NOR2B
      port map(A => N_22_0_0, B => \data_counter[7]_net_1\, Y => 
        N_23_0_0);
    
    \state_RNI6D91[2]\ : OR2
      port map(A => \state[4]_net_1\, B => \state[2]_net_1\, Y
         => N_518_1);
    
    \data_counter[3]\ : DFN1C0
      port map(D => N_192, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_counter[3]_net_1\);
    
    \DMAIn.Address_RNI9IRJ[23]\ : MX2
      port map(A => \Address[23]\, B => data_address(23), S => 
        time_select_0, Y => N_970);
    
    \state[5]\ : DFN1P0
      port map(D => N_4, CLK => HCLK_c, PRE => HRESETn_c, Q => 
        \state[5]_net_1\);
    
    \grant_counter_RNO[30]\ : XA1
      port map(A => \grant_counter[30]_net_1\, B => I129_un1_Y, C
         => N_202, Y => N_141);
    
    \data_counter_RNO[8]\ : XA1B
      port map(A => \data_counter[8]_net_1\, B => N_23_0_0, C => 
        N_198_0, Y => \data_counter_8[8]\);
    
    \data_counter[28]\ : DFN1C0
      port map(D => \data_counter_8[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[28]_net_1\);
    
    \state_RNI9EI2[0]\ : OR2
      port map(A => N_518_1, B => N_338_1, Y => N_516);
    
    \data_counter[10]\ : DFN1C0
      port map(D => \data_counter_8[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[10]_net_1\);
    
    \data_counter_RNO[13]\ : XA1C
      port map(A => \data_counter[13]_net_1\, B => N_28_0, C => 
        N_198_0, Y => \data_counter_8[13]\);
    
    \data_counter[12]\ : DFN1C0
      port map(D => \data_counter_8[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[12]_net_1\);
    
    \data_counter[24]\ : DFN1C0
      port map(D => \data_counter_8[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[24]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DMAIn.Address_RNO[26]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(26), Y
         => N_71);
    
    un1_state_4_m23 : NOR2B
      port map(A => N_23_0_0, B => \data_counter[8]_net_1\, Y => 
        N_24_0_0);
    
    un1_hresetn_inv_2_m47 : NOR3C
      port map(A => \grant_counter[15]_net_1\, B => N_44, C => 
        \grant_counter[16]_net_1\, Y => N_48);
    
    \DMAIn.Address_RNO[23]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(23), Y
         => N_65);
    
    \DMAIn.Address_RNIOUQJ[19]\ : MX2
      port map(A => \Address[19]\, B => data_address(19), S => 
        time_select_0, Y => N_966);
    
    \DMAIn.Address[12]\ : DFN1E1C0
      port map(D => N_43, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[12]\);
    
    \data_counter_RNIQ8473[22]\ : NOR3C
      port map(A => un1_state_5_i_o2_21, B => un1_state_5_i_o2_20, 
        C => un1_state_5_i_o2_27, Y => un1_state_5_i_o2_29);
    
    \data_counter[27]\ : DFN1C0
      port map(D => \data_counter_8[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[27]_net_1\);
    
    \grant_counter_RNO[1]\ : AO1
      port map(A => N_31_0_i_0, B => N_202, C => N_513, Y => 
        \grant_counter_RNO[1]_net_1\);
    
    \DMAIn.Address[5]\ : DFN1E1C0
      port map(D => N_23, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[5]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \data_counter_RNO[10]\ : XA1B
      port map(A => \data_counter[10]_net_1\, B => N_25_0_0, C
         => N_198_0, Y => \data_counter_8[10]\);
    
    \data_counter_RNICTS71[2]\ : NOR3C
      port map(A => un1_state_5_i_o2_13, B => un1_state_5_i_o2_12, 
        C => un1_state_5_i_o2_23, Y => un1_state_5_i_o2_27);
    
    \grant_counter_RNO[28]\ : NOR2A
      port map(A => N_202, B => \un1_hresetn_inv_2_i[3]\, Y => 
        N_137);
    
    \grant_counter[17]\ : DFN1
      port map(D => N_115, CLK => HCLK_c, Q => 
        \grant_counter[17]_net_1\);
    
    \grant_counter_RNINSC[16]\ : NOR2
      port map(A => \grant_counter[16]_net_1\, B => 
        \grant_counter[17]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_9[3]\);
    
    \data_counter_RNO[27]\ : XA1B
      port map(A => \data_counter[27]_net_1\, B => N_68_0, C => 
        N_198, Y => \data_counter_8[27]\);
    
    \grant_counter_RNO[24]\ : NOR2A
      port map(A => N_202, B => \un1_hresetn_inv_2_i[7]\, Y => 
        N_129);
    
    \data_counter[1]\ : DFN1C0
      port map(D => N_188, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_counter[1]_net_1\);
    
    \grant_counter_RNO[10]\ : XA1
      port map(A => \grant_counter[10]_net_1\, B => N_25_0, C => 
        N_202_0, Y => N_101);
    
    \grant_counter[30]\ : DFN1
      port map(D => N_141, CLK => HCLK_c, Q => 
        \grant_counter[30]_net_1\);
    
    \grant_counter[9]\ : DFN1
      port map(D => N_99, CLK => HCLK_c, Q => 
        \grant_counter[9]_net_1\);
    
    \data_counter_RNO_1[0]\ : NOR3
      port map(A => N_235, B => \state[0]_net_1\, C => N_508, Y
         => N_339);
    
    \data_counter_RNO[6]\ : XA1B
      port map(A => \data_counter[6]_net_1\, B => N_21_0_0, C => 
        N_198, Y => \data_counter_8[6]\);
    
    \state_RNI1BT21[3]\ : OR2A
      port map(A => N_348, B => \state[3]_net_1\, Y => N_509);
    
    \DMAIn.Address_RNO[30]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(30), Y
         => N_79);
    
    \grant_counter_RNIFSC[12]\ : NOR2
      port map(A => \grant_counter[12]_net_1\, B => 
        \grant_counter[13]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_7[3]\);
    
    un1_state_4_m57 : NOR2B
      port map(A => N_56_0, B => \data_counter[21]_net_1\, Y => 
        N_58);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_7 : NOR2B
      port map(A => \grant_counter[28]_net_1\, B => 
        \grant_counter[29]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_7);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_4 : NOR2B
      port map(A => \grant_counter[22]_net_1\, B => 
        \grant_counter[23]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_4);
    
    \grant_counter_RNO[12]\ : XA1
      port map(A => \grant_counter[12]_net_1\, B => N_27_0, C => 
        N_202_0, Y => N_105);
    
    \DMAIn.Address_RNO[8]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(8), Y
         => N_29);
    
    \DMAIn.Address[9]\ : DFN1E1C0
      port map(D => N_31, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[9]\);
    
    un1_state_4_m61 : NOR2B
      port map(A => N_60_0, B => \data_counter[23]_net_1\, Y => 
        N_62);
    
    un1_state_4_m26 : OR2B
      port map(A => N_26_0_0, B => \data_counter[11]_net_1\, Y
         => N_27_0_0);
    
    \grant_counter[18]\ : DFN1
      port map(D => N_117, CLK => HCLK_c, Q => 
        \grant_counter[18]_net_1\);
    
    \data_counter_RNO[4]\ : XA1B
      port map(A => \data_counter[4]_net_1\, B => N_19_0_0, C => 
        N_198, Y => \data_counter_8[4]\);
    
    \data_counter[29]\ : DFN1C0
      port map(D => \data_counter_8[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[29]_net_1\);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_1 : NOR2B
      port map(A => \grant_counter[16]_net_1\, B => 
        \grant_counter[17]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_1);
    
    \DMAIn.Address_RNO[18]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(18), Y
         => N_55);
    
    \DMAIn.Address[10]\ : DFN1E1C0
      port map(D => N_33, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[10]\);
    
    un1_state_4_m31 : AX1E
      port map(A => \data_counter[1]_net_1\, B => N_16_0, C => 
        \data_counter[2]_net_1\, Y => \un1_state_4_i[29]\);
    
    \DMAIn.Address_RNO[29]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(29), Y
         => N_77);
    
    \state_RNI1E9S2[3]\ : OAI1
      port map(A => N_246, B => un1_state_7_i_a4_0_1, C => N_516, 
        Y => N_146);
    
    un1_state_4_m32 : XNOR2
      port map(A => N_18_0, B => \data_counter[3]_net_1\, Y => 
        \un1_state_4_i[28]\);
    
    \DMAIn.Address_RNID6SJ[31]\ : MX2
      port map(A => \Address[31]\, B => data_address(31), S => 
        time_select_0, Y => N_978);
    
    \data_counter[2]\ : DFN1C0
      port map(D => N_190, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_counter[2]_net_1\);
    
    un1_hresetn_inv_2_m67 : NOR3C
      port map(A => \grant_counter[25]_net_1\, B => N_64, C => 
        \grant_counter[26]_net_1\, Y => N_68);
    
    un1_hresetn_inv_2_m43_m6_0_a2_2 : NOR2B
      port map(A => \grant_counter[10]_net_1\, B => 
        \grant_counter[11]_net_1\, Y => m43_m6_0_a2_2);
    
    \DMAIn.Address_RNI86SJ[30]\ : MX2
      port map(A => \Address[30]\, B => data_address(30), S => 
        time_select_0, Y => N_977);
    
    \DMAIn.Address[11]\ : DFN1E1C0
      port map(D => N_35, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[11]\);
    
    un1_hresetn_inv_2_m34 : AX1E
      port map(A => \grant_counter[4]_net_1\, B => N_19_0, C => 
        \grant_counter[5]_net_1\, Y => \un1_hresetn_inv_2_i[26]\);
    
    \state_RNIR8B01[4]\ : OR2B
      port map(A => \state[4]_net_1\, B => Grant, Y => \N_200\);
    
    \grant_counter[21]\ : DFN1
      port map(D => N_123, CLK => HCLK_c, Q => 
        \grant_counter[21]_net_1\);
    
    \DMAIn.Address_RNI6EA51[9]\ : MX2
      port map(A => \Address[9]\, B => data_address(9), S => 
        time_select, Y => N_956);
    
    \DMAIn.Address_RNI2JRJ[28]\ : MX2C
      port map(A => \Address[28]\, B => data_address(28), S => 
        time_select_0, Y => N_975);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_7 : NOR2B
      port map(A => \data_counter[28]_net_1\, B => 
        \data_counter[29]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_7_0);
    
    \grant_counter[22]\ : DFN1
      port map(D => N_125, CLK => HCLK_c, Q => 
        \grant_counter[22]_net_1\);
    
    \DMAIn.Address[14]\ : DFN1E1C0
      port map(D => N_47, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[14]\);
    
    \DMAIn.Burst_RNI9478\ : OR2A
      port map(A => Burst, B => time_select, Y => un7_dmain(66));
    
    un1_state_4_m63 : NOR2B
      port map(A => N_62, B => \data_counter[24]_net_1\, Y => 
        N_64_0);
    
    un1_state_4_m44 : AX1E
      port map(A => \data_counter[14]_net_1\, B => N623_0, C => 
        \data_counter[15]_net_1\, Y => N_45);
    
    \state_RNISRSN8[3]\ : OR2B
      port map(A => N_509, B => N_344, Y => N_198);
    
    \DMAIn.Address_RNITB461[8]\ : MX2
      port map(A => \Address[8]\, B => data_address(8), S => 
        time_select, Y => N_955);
    
    \state_RNO_0[0]\ : NOR2A
      port map(A => \state[0]_net_1\, B => Ready, Y => 
        \state_RNO_0[0]_net_1\);
    
    \grant_counter_RNO[18]\ : NOR2A
      port map(A => N_202_0, B => \un1_hresetn_inv_2_i[13]\, Y
         => N_117);
    
    \data_counter[0]\ : DFN1C0
      port map(D => N_186, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_counter[0]_net_1\);
    
    un1_hresetn_inv_2_m51 : NOR3C
      port map(A => \grant_counter[17]_net_1\, B => N_48, C => 
        \grant_counter[18]_net_1\, Y => N_52);
    
    \grant_counter_RNO[27]\ : XA1
      port map(A => \grant_counter[27]_net_1\, B => N_68, C => 
        N_202, Y => N_135);
    
    \DMAIn.Address_RNO[16]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(16), Y
         => N_51);
    
    \grant_counter_RNO[14]\ : XA1
      port map(A => \grant_counter[14]_net_1\, B => N623, C => 
        N_202_0, Y => N_109);
    
    un1_state_4_m59 : NOR2B
      port map(A => N_58, B => \data_counter[22]_net_1\, Y => 
        N_60_0);
    
    \data_counter_RNI1O34[8]\ : NOR2
      port map(A => \data_counter[8]_net_1\, B => 
        \data_counter[9]_net_1\, Y => un1_state_5_i_o2_4);
    
    un1_hresetn_inv_2_m50 : AX1E
      port map(A => \grant_counter[17]_net_1\, B => N_48, C => 
        \grant_counter[18]_net_1\, Y => \un1_hresetn_inv_2_i[13]\);
    
    \DMAIn.Address_RNO[13]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(13), Y
         => N_45_0);
    
    un1_state_4_m25 : NOR2B
      port map(A => N_25_0_0, B => \data_counter[10]_net_1\, Y
         => N_26_0_0);
    
    \grant_counter_RNIU9Q[26]\ : NOR3A
      port map(A => \state_ns_i_a2_0_i_o2_15[3]\, B => 
        \grant_counter[27]_net_1\, C => \grant_counter[26]_net_1\, 
        Y => \state_ns_i_a2_0_i_o2_23[3]\);
    
    \DMAIn.Address_RNIKHKI[10]\ : MX2
      port map(A => \Address[10]\, B => data_address(10), S => 
        time_select, Y => N_957);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state_RNIS4Q9[3]\ : OR3A
      port map(A => Ready, B => \state[3]_net_1\, C => N_518_1, Y
         => un1_state_7_i_a4_0_1);
    
    \DMAIn.Address_RNO[7]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(7), Y
         => N_27);
    
    \data_counter_RNO_2[0]\ : NOR3B
      port map(A => N_235, B => \state[3]_net_1\, C => 
        \un1_state_4_i_i[31]\, Y => N_336);
    
    \data_counter_RNO[16]\ : XA1B
      port map(A => \data_counter[16]_net_1\, B => N_46, C => 
        N_198_0, Y => \data_counter_8[16]\);
    
    \data_counter_RNO[29]\ : XA1B
      port map(A => \data_counter[29]_net_1\, B => N_72_0, C => 
        N_198, Y => \data_counter_8[29]\);
    
    un1_hresetn_inv_2_m16 : NOR3C
      port map(A => \grant_counter[0]_net_1\, B => 
        un1_hresetn_inv_i_0, C => \grant_counter[1]_net_1\, Y => 
        N_17_0);
    
    \DMAIn.Address[8]\ : DFN1E1C0
      port map(D => N_29, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[8]\);
    
    \state_RNO[4]\ : AO1A
      port map(A => Grant, B => \state[4]_net_1\, C => Request_5, 
        Y => N_84);
    
    \state_RNIK8SG_0[3]\ : OR2A
      port map(A => \state[3]_net_1\, B => Fault, Y => N_522);
    
    un1_state_4_m27_m6_0_a2 : OR2B
      port map(A => m27_m6_0_a2_4, B => N_19_0_0, Y => N_28_0);
    
    \grant_counter_RNIP4D[24]\ : NOR2
      port map(A => \grant_counter[24]_net_1\, B => 
        \grant_counter[25]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_13[3]\);
    
    \state_RNIAMD44[4]\ : NOR3A
      port map(A => un1_hresetn_inv_i_0, B => N_246, C => 
        \state[4]_net_1\, Y => N_513);
    
    \DMAIn.Address_RNO[19]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(19), Y
         => N_57);
    
    \DMAIn.Address[0]\ : DFN1E1C0
      port map(D => N_13, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[0]\);
    
    un1_hresetn_inv_2_m25 : NOR2B
      port map(A => N_25_0, B => \grant_counter[10]_net_1\, Y => 
        N_26_0);
    
    un1_state_4_m27_m6_0_a2_4_5 : NOR3C
      port map(A => \data_counter[6]_net_1\, B => 
        \data_counter[5]_net_1\, C => m27_m6_0_a2_4_2, Y => 
        m27_m6_0_a2_4_5);
    
    \state_RNO[2]\ : AO1C
      port map(A => N_346, B => N_246, C => N_522, Y => N_151);
    
    \grant_counter_RNO[17]\ : XA1
      port map(A => \grant_counter[17]_net_1\, B => N_48, C => 
        N_202_0, Y => N_115);
    
    \grant_counter_RNIM2O7[30]\ : NOR2
      port map(A => \grant_counter[5]_net_1\, B => 
        \grant_counter[30]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_1[3]\);
    
    \state_RNIQIK31[4]\ : OR2A
      port map(A => HRESETn_c, B => \N_200\, Y => N_202);
    
    un1_state_4_m71 : NOR2B
      port map(A => N_70, B => \data_counter[28]_net_1\, Y => 
        N_72_0);
    
    \grant_counter[10]\ : DFN1
      port map(D => N_101, CLK => HCLK_c, Q => 
        \grant_counter[10]_net_1\);
    
    \data_counter_RNO[28]\ : XA1B
      port map(A => \data_counter[28]_net_1\, B => N_70, C => 
        N_198, Y => \data_counter_8[28]\);
    
    \grant_counter[24]\ : DFN1
      port map(D => N_129, CLK => HCLK_c, Q => 
        \grant_counter[24]_net_1\);
    
    \data_counter_RNO[15]\ : NOR2
      port map(A => N_45, B => N_198_0, Y => \data_counter_8[15]\);
    
    \DMAIn.Lock_RNILJE7\ : MX2C
      port map(A => Lock, B => Lock_0, S => time_select, Y => 
        N_1013);
    
    un1_state_4_m65 : NOR2B
      port map(A => N_64_0, B => \data_counter[25]_net_1\, Y => 
        N_66);
    
    \DMAIn.Address_RNI4IRJ[22]\ : MX2
      port map(A => \Address[22]\, B => data_address(22), S => 
        time_select_0, Y => N_969);
    
    \grant_counter[16]\ : DFN1
      port map(D => N_113, CLK => HCLK_c, Q => 
        \grant_counter[16]_net_1\);
    
    \DMAIn.Address_RNION361[7]\ : MX2
      port map(A => \Address[7]\, B => data_address(7), S => 
        time_select, Y => N_954);
    
    \DMAIn.Address[15]\ : DFN1E1C0
      port map(D => N_49, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[15]\);
    
    un1_state_4_m20 : NOR2B
      port map(A => N_20_0, B => \data_counter[5]_net_1\, Y => 
        N_21_0_0);
    
    \state_RNIAC4L7[3]\ : AO1D
      port map(A => N_241, B => N_235, C => N_242, Y => N_154);
    
    \grant_counter[19]\ : DFN1
      port map(D => N_119, CLK => HCLK_c, Q => 
        \grant_counter[19]_net_1\);
    
    send_ok_RNIC0Q : NOR2
      port map(A => data_send_ok, B => data_send_ko, Y => 
        un1_data_send_ok);
    
    un1_hresetn_inv_2_m32 : AX1C
      port map(A => \grant_counter[2]_net_1\, B => N_17_0, C => 
        \grant_counter[3]_net_1\, Y => N_33_0_i_0);
    
    un1_hresetn_inv_2_m27 : NOR2B
      port map(A => N_27_0, B => \grant_counter[12]_net_1\, Y => 
        N_28_0_0);
    
    \data_counter[18]\ : DFN1C0
      port map(D => \data_counter_8[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[18]_net_1\);
    
    \DMAIn.Address_RNO[3]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(3), Y
         => N_19);
    
    \data_counter_RNO[24]\ : XA1B
      port map(A => \data_counter[24]_net_1\, B => N_62, C => 
        N_198, Y => \data_counter_8[24]\);
    
    \data_counter[14]\ : DFN1C0
      port map(D => \data_counter_8[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[14]_net_1\);
    
    \grant_counter_RNO[23]\ : XA1
      port map(A => \grant_counter[23]_net_1\, B => N_60, C => 
        N_202, Y => N_127);
    
    \DMAIn.Address_RNI5TN41[3]\ : MX2
      port map(A => \Address[3]\, B => data_address(3), S => 
        time_select_0, Y => N_950);
    
    un1_state_4_m28_m6_0 : NOR2B
      port map(A => \data_counter[13]_net_1\, B => 
        \data_counter[1]_net_1\, Y => m28_m6_0);
    
    \state_RNIK8SG[3]\ : OR2B
      port map(A => \state[3]_net_1\, B => Fault, Y => N_241);
    
    \DMAIn.Request_RNIJKMF\ : MX2
      port map(A => Request, B => Request_0, S => time_select, Y
         => N_1011);
    
    \DMAIn.Address_RNO[21]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(21), Y
         => N_61);
    
    \DMAIn.Address[23]\ : DFN1E1C0
      port map(D => N_65, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[23]\);
    
    \grant_counter[23]\ : DFN1
      port map(D => N_127, CLK => HCLK_c, Q => 
        \grant_counter[23]_net_1\);
    
    \data_counter[17]\ : DFN1C0
      port map(D => \data_counter_8[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[17]_net_1\);
    
    \state_RNIAC4L7_0[3]\ : AO1D
      port map(A => N_241, B => N_235, C => N_242, Y => N_154_0);
    
    \state_RNI3191[1]\ : NOR2
      port map(A => \state[1]_net_1\, B => \state[2]_net_1\, Y
         => un1_state_2_i_o2_0);
    
    \grant_counter_RNIH4D[20]\ : NOR2
      port map(A => \grant_counter[20]_net_1\, B => 
        \grant_counter[21]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_11[3]\);
    
    \DMAIn.Address_RNIQKM41[1]\ : MX2
      port map(A => \Address[1]\, B => data_address(1), S => 
        time_select_0, Y => N_948);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_14 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_9_0, B => 
        ADD_32x32_fast_I129_un1_Y_8_0, C => 
        ADD_32x32_fast_I129_un1_Y_13_0, Y => 
        ADD_32x32_fast_I129_un1_Y_14_0);
    
    \data_counter_RNIJN34[3]\ : NOR2B
      port map(A => \data_counter[3]_net_1\, B => 
        \data_counter[0]_net_1\, Y => un1_state_5_i_o2_15);
    
    \data_counter[31]\ : DFN1C0
      port map(D => \data_counter_8[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[31]_net_1\);
    
    \data_counter_RNILUOF[20]\ : NOR2
      port map(A => \data_counter[20]_net_1\, B => 
        \data_counter[21]_net_1\, Y => un1_state_5_i_o2_9);
    
    un1_state_4_m29 : XNOR2
      port map(A => \data_counter[0]_net_1\, B => N_510, Y => 
        \un1_state_4_i_i[31]\);
    
    un1_hresetn_inv_2_m28 : NOR2B
      port map(A => N_28_0_0, B => \grant_counter[13]_net_1\, Y
         => N623);
    
    \data_counter_RNO_0[0]\ : AO1D
      port map(A => N_508, B => N_338_1, C => N_337, Y => 
        \data_counter_8_i_0[0]\);
    
    \data_counter_RNIOTJV[18]\ : NOR3A
      port map(A => un1_state_5_i_o2_9, B => 
        \data_counter[19]_net_1\, C => \data_counter[18]_net_1\, 
        Y => un1_state_5_i_o2_20);
    
    \grant_counter[31]\ : DFN1
      port map(D => N_143, CLK => HCLK_c, Q => 
        \grant_counter[31]_net_1\);
    
    \grant_counter[15]\ : DFN1
      port map(D => N_111, CLK => HCLK_c, Q => 
        \grant_counter[15]_net_1\);
    
    \DMAIn.Address_RNO[1]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(1), Y
         => N_15);
    
    \grant_counter[6]\ : DFN1
      port map(D => N_93, CLK => HCLK_c, Q => 
        \grant_counter[6]_net_1\);
    
    \DMAIn.Address_RNO[22]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(22), Y
         => N_63);
    
    \data_counter[19]\ : DFN1C0
      port map(D => \data_counter_8[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[19]_net_1\);
    
    \DMAIn.Address[16]\ : DFN1E1C0
      port map(D => N_51, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[16]\);
    
    \grant_counter_RNO_0[0]\ : XA1A
      port map(A => \grant_counter[0]_net_1\, B => 
        un1_hresetn_inv_i_0, C => N_202_0, Y => 
        \grant_counter_0_0_0[0]\);
    
    \grant_counter[8]\ : DFN1
      port map(D => N_97, CLK => HCLK_c, Q => 
        \grant_counter[8]_net_1\);
    
    \data_counter_RNIN6PF[30]\ : NOR2
      port map(A => \data_counter[13]_net_1\, B => 
        \data_counter[30]_net_1\, Y => un1_state_5_i_o2_1);
    
    \state_RNI3191[0]\ : OR2
      port map(A => \state[3]_net_1\, B => \state[0]_net_1\, Y
         => N_338_1);
    
    un1_state_4_m30 : XNOR2
      port map(A => N_16_0, B => \data_counter[1]_net_1\, Y => 
        \un1_state_4_i[30]\);
    
    \DMAIn.Address_RNO[24]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(24), Y
         => N_67);
    
    \data_counter_RNO[3]\ : AOI1B
      port map(A => \un1_state_4_i[28]\, B => N_344, C => N_509, 
        Y => N_192);
    
    un1_hresetn_inv_2_m43_m6_0_a2_5 : NOR3C
      port map(A => \grant_counter[9]_net_1\, B => 
        \grant_counter[8]_net_1\, C => m43_m6_0_a2_2, Y => 
        m43_m6_0_a2_5);
    
    \DMAIn.Address_RNO[25]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(25), Y
         => N_69);
    
    \data_counter_RNO[5]\ : XA1B
      port map(A => \data_counter[5]_net_1\, B => N_20_0, C => 
        N_198, Y => \data_counter_8[5]\);
    
    \data_counter_RNITUPF[24]\ : NOR2
      port map(A => \data_counter[24]_net_1\, B => 
        \data_counter[25]_net_1\, Y => un1_state_5_i_o2_11);
    
    un1_state_4_m67 : NOR2B
      port map(A => N_66, B => \data_counter[26]_net_1\, Y => 
        N_68_0);
    
    \grant_counter_RNO[13]\ : XA1
      port map(A => \grant_counter[13]_net_1\, B => N_28_0_0, C
         => N_202_0, Y => N_107);
    
    \grant_counter_RNIDK1F[1]\ : NOR2B
      port map(A => \grant_counter[0]_net_1\, B => 
        \grant_counter[1]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_2[3]\);
    
    \state[3]\ : DFN1C0
      port map(D => \state_RNO[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    
    \state_RNIJKJ6[1]\ : AO1A
      port map(A => data_send, B => \state_0[5]_net_1\, C => 
        \state[1]_net_1\, Y => \state_ns_i_a2_i_0_0[0]\);
    
    \data_counter[7]\ : DFN1C0
      port map(D => \data_counter_8[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[7]_net_1\);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_14 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_9, B => 
        ADD_32x32_fast_I129_un1_Y_8, C => 
        ADD_32x32_fast_I129_un1_Y_13, Y => 
        ADD_32x32_fast_I129_un1_Y_14);
    
    \grant_counter_RNO[21]\ : XA1
      port map(A => \grant_counter[21]_net_1\, B => N_56, C => 
        N_202, Y => N_123);
    
    \data_counter[5]\ : DFN1C0
      port map(D => \data_counter_8[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[5]_net_1\);
    
    \DMAIn.Request\ : DFN1E1C0
      port map(D => Request_5, CLK => HCLK_c, CLR => HRESETn_c, E
         => N_156, Q => Request);
    
    \DMAIn.Address_RNO[11]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(11), Y
         => N_35);
    
    \grant_counter_RNO_0[4]\ : AO1C
      port map(A => N_246, B => un1_hresetn_inv_i_0, C => N_202_0, 
        Y => \grant_counter_0_i_0[4]\);
    
    \DMAIn.Address_RNO[6]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(6), Y
         => N_25);
    
    \DMAIn.Address[17]\ : DFN1E1C0
      port map(D => N_53, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[17]\);
    
    \data_counter_RNIVEQF[16]\ : NOR2
      port map(A => \data_counter[16]_net_1\, B => 
        \data_counter[17]_net_1\, Y => un1_state_5_i_o2_7);
    
    \grant_counter_RNO[31]\ : XA1
      port map(A => \grant_counter[31]_net_1\, B => N_75, C => 
        N_202, Y => N_143);
    
    \grant_counter_RNIGI0V[6]\ : NOR3C
      port map(A => \state_ns_i_a2_0_i_o2_5[3]\, B => 
        \state_ns_i_a2_0_i_o2_4[3]\, C => 
        \state_ns_i_a2_0_i_o2_19[3]\, Y => 
        \state_ns_i_a2_0_i_o2_25[3]\);
    
    \state_RNIEK821[0]\ : NOR2
      port map(A => \state[0]_net_1\, B => N_243, Y => N_348);
    
    un1_state_4_m28_m6_5 : AOI1B
      port map(A => \state[3]_net_1\, B => OKAY, C => m28_m6_4, Y
         => m28_m6_5);
    
    \state_RNIF6GI1[0]\ : OR2A
      port map(A => N_348, B => OKAY, Y => N_510);
    
    \DMAIn.Address[22]\ : DFN1E1C0
      port map(D => N_63, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[22]\);
    
    \data_counter_RNO[30]\ : NOR2
      port map(A => \un1_state_4_i[1]\, B => N_198, Y => 
        \data_counter_8[30]\);
    
    \data_counter[9]\ : DFN1C0
      port map(D => \data_counter_8[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[9]_net_1\);
    
    un1_state_4_m69 : NOR2B
      port map(A => N_68_0, B => \data_counter[27]_net_1\, Y => 
        N_70);
    
    un1_hresetn_inv_2_m43_m6_0_a2_4 : NOR3C
      port map(A => \grant_counter[7]_net_1\, B => 
        \grant_counter[6]_net_1\, C => \grant_counter[14]_net_1\, 
        Y => m43_m6_0_a2_4);
    
    un1_state_4_m27_m6_0_a2_4 : NOR3C
      port map(A => m27_m6_0_a2_4_4, B => m27_m6_0_a2_4_3, C => 
        m27_m6_0_a2_4_5, Y => m27_m6_0_a2_4);
    
    \data_counter[30]\ : DFN1C0
      port map(D => \data_counter_8[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[30]_net_1\);
    
    un1_state_4_m28_m6_1 : NOR2B
      port map(A => \data_counter[2]_net_1\, B => 
        \data_counter[3]_net_1\, Y => m28_m6_1);
    
    \data_counter_RNO[7]\ : XA1B
      port map(A => \data_counter[7]_net_1\, B => N_22_0_0, C => 
        N_198_0, Y => \data_counter_8[7]\);
    
    \data_counter_RNO[11]\ : XA1B
      port map(A => \data_counter[11]_net_1\, B => N_26_0_0, C
         => N_198_0, Y => \data_counter_8[11]\);
    
    un1_hresetn_inv_2_m62 : AX1E
      port map(A => \grant_counter[23]_net_1\, B => N_60, C => 
        \grant_counter[24]_net_1\, Y => \un1_hresetn_inv_2_i[7]\);
    
    \grant_counter_RNO[2]\ : AO1
      port map(A => N_32_0_i_0, B => N_202, C => N_513, Y => 
        \grant_counter_RNO[2]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \data_counter_RNO[23]\ : XA1B
      port map(A => \data_counter[23]_net_1\, B => N_60_0, C => 
        N_198, Y => \data_counter_8[23]\);
    
    un1_hresetn_inv_2_m24 : NOR2B
      port map(A => N_24_0, B => \grant_counter[9]_net_1\, Y => 
        N_25_0);
    
    \DMAIn.Address_RNO[12]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(12), Y
         => N_43);
    
    un1_hresetn_inv_2_m55 : NOR3C
      port map(A => \grant_counter[19]_net_1\, B => N_52, C => 
        \grant_counter[20]_net_1\, Y => N_56);
    
    \grant_counter_RNO[25]\ : XA1
      port map(A => \grant_counter[25]_net_1\, B => N_64, C => 
        N_202, Y => N_131);
    
    \DMAIn.Address_RNITIRJ[27]\ : MX2C
      port map(A => \Address[27]\, B => data_address(27), S => 
        time_select_0, Y => N_974);
    
    \DMAIn.Address_RNO[14]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(14), Y
         => N_47);
    
    \grant_counter_RNO[11]\ : XA1
      port map(A => \grant_counter[11]_net_1\, B => N_26_0, C => 
        N_202_0, Y => N_103);
    
    \grant_counter_RNI2E83[14]\ : NOR3C
      port map(A => \state_ns_i_a2_0_i_o2_21[3]\, B => 
        \state_ns_i_a2_0_i_o2_20[3]\, C => 
        \state_ns_i_a2_0_i_o2_27[3]\, Y => 
        \state_ns_i_a2_0_i_o2_29[3]\);
    
    \DMAIn.Address[20]\ : DFN1E1C0
      port map(D => N_59, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[20]\);
    
    \DMAIn.Address_RNO[15]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(15), Y
         => N_49);
    
    un1_state_4_m74_0 : NOR2B
      port map(A => \data_counter[30]_net_1\, B => 
        \data_counter[29]_net_1\, Y => m74_0);
    
    \DMAIn.Address_RNIOIRJ[26]\ : MX2C
      port map(A => \Address[26]\, B => data_address(26), S => 
        time_select_0, Y => N_973);
    
    \data_counter_RNO[20]\ : XA1B
      port map(A => \data_counter[20]_net_1\, B => N_54, C => 
        N_198_0, Y => \data_counter_8[20]\);
    
    \state_RNI2R0V2[1]\ : AO1D
      port map(A => N_346, B => N_246, C => 
        \state_ns_i_a2_i_0_0[0]\, Y => N_4);
    
    \DMAIn.Address_RNI7JRJ[29]\ : MX2
      port map(A => \Address[29]\, B => data_address(29), S => 
        time_select_0, Y => N_976);
    
    \DMAIn.Address[21]\ : DFN1E1C0
      port map(D => N_61, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[21]\);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_13 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_5_0, B => 
        ADD_32x32_fast_I129_un1_Y_4_0, C => 
        ADD_32x32_fast_I129_un1_Y_11_0, Y => 
        ADD_32x32_fast_I129_un1_Y_13_0);
    
    \grant_counter[5]\ : DFN1
      port map(D => N_91, CLK => HCLK_c, Q => 
        \grant_counter[5]_net_1\);
    
    \DMAIn.Address_RNO[9]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(9), Y
         => N_31);
    
    \DMAIn.Address[18]\ : DFN1E1C0
      port map(D => N_55, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[18]\);
    
    \data_counter[25]\ : DFN1C0
      port map(D => \data_counter_8[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[25]_net_1\);
    
    \grant_counter[4]\ : DFN1
      port map(D => N_89, CLK => HCLK_c, Q => 
        \grant_counter[4]_net_1\);
    
    \grant_counter[11]\ : DFN1
      port map(D => N_103, CLK => HCLK_c, Q => 
        \grant_counter[11]_net_1\);
    
    \DMAIn.Address[24]\ : DFN1E1C0
      port map(D => N_67, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[24]\);
    
    \grant_counter[12]\ : DFN1
      port map(D => N_105, CLK => HCLK_c, Q => 
        \grant_counter[12]_net_1\);
    
    \DMAIn.Burst_RNO\ : NOR3C
      port map(A => N_522, B => Burst, C => N_526, Y => N_194_i_0);
    
    un1_hresetn_inv_2_m43_m6_0_a2 : NOR3C
      port map(A => m43_m6_0_a2_6, B => m43_m6_0_a2_5, C => 
        N_21_0, Y => N_44);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_9 : NOR3C
      port map(A => \grant_counter[19]_net_1\, B => 
        \grant_counter[18]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_3, Y => 
        ADD_32x32_fast_I129_un1_Y_9);
    
    \DMAIn.Address[19]\ : DFN1E1C0
      port map(D => N_57, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154_0, Q => \Address[19]\);
    
    \data_counter_RNO[1]\ : AOI1B
      port map(A => \un1_state_4_i[30]\, B => N_344, C => N_509, 
        Y => N_188);
    
    \state_RNIMV7G3[3]\ : OR3B
      port map(A => \state[3]_net_1\, B => Grant, C => N_246, Y
         => N_526);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_4 : NOR2B
      port map(A => \data_counter[22]_net_1\, B => 
        \data_counter[23]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_4_0);
    
    \state_RNISRSN8_0[3]\ : OR2B
      port map(A => N_509, B => N_344, Y => N_198_0);
    
    un1_hresetn_inv_2_m74 : NOR3C
      port map(A => \grant_counter[29]_net_1\, B => 
        \grant_counter[30]_net_1\, C => N_72, Y => N_75);
    
    \grant_counter_RNI15D[28]\ : NOR2
      port map(A => \grant_counter[28]_net_1\, B => 
        \grant_counter[29]_net_1\, Y => 
        \state_ns_i_a2_0_i_o2_15[3]\);
    
    \data_counter[4]\ : DFN1C0
      port map(D => \data_counter_8[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[4]_net_1\);
    
    \DMAIn.Address_RNIVHRJ[21]\ : MX2
      port map(A => \Address[21]\, B => data_address(21), S => 
        time_select_0, Y => N_968);
    
    \grant_counter_RNO[15]\ : XA1
      port map(A => \grant_counter[15]_net_1\, B => N_44, C => 
        N_202_0, Y => N_111);
    
    un1_hresetn_inv_2_m43_m6_0_a2_6 : NOR3C
      port map(A => \grant_counter[13]_net_1\, B => 
        \grant_counter[12]_net_1\, C => m43_m6_0_a2_4, Y => 
        m43_m6_0_a2_6);
    
    \grant_counter[7]\ : DFN1
      port map(D => N_95, CLK => HCLK_c, Q => 
        \grant_counter[7]_net_1\);
    
    \DMAIn.Address_RNO[31]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_address(31), Y
         => N_81);
    
    \state[2]\ : DFN1C0
      port map(D => N_151, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[2]_net_1\);
    
    \data_counter_RNIE4HJ1[8]\ : NOR3C
      port map(A => un1_state_5_i_o2_5, B => un1_state_5_i_o2_4, 
        C => un1_state_5_i_o2_19, Y => un1_state_5_i_o2_25);
    
    send_ko : DFN1E1C0
      port map(D => \state[1]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_146, Q => data_send_ko);
    
    \data_counter_RNO[12]\ : XA1C
      port map(A => \data_counter[12]_net_1\, B => N_27_0_0, C
         => N_198_0, Y => \data_counter_8[12]\);
    
    un1_state_4_ADD_32x32_fast_I190_Y_0 : AX1E
      port map(A => N623_0, B => ADD_32x32_fast_I129_un1_Y_14_0, 
        C => \data_counter[30]_net_1\, Y => \un1_state_4_i[1]\);
    
    \DMAIn.Address_RNIMC0J[18]\ : MX2
      port map(A => \Address[18]\, B => data_address(18), S => 
        time_select_0, Y => N_965);
    
    un1_hresetn_inv_2_m31 : XOR2
      port map(A => N_17_0, B => \grant_counter[2]_net_1\, Y => 
        N_32_0_i_0);
    
    un1_state_4_m27_m6_0_a2_4_3 : NOR2B
      port map(A => \data_counter[9]_net_1\, B => 
        \data_counter[10]_net_1\, Y => m27_m6_0_a2_4_3);
    
    \DMAIn.Store\ : DFN1E1C0
      port map(D => \state[5]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_156, Q => Store);
    
    \DMAIn.Address_RNI9R161[4]\ : MX2
      port map(A => \Address[4]\, B => data_address(4), S => 
        time_select, Y => N_951);
    
    un1_state_4_m27_m6_0_a2_4_2 : NOR2B
      port map(A => \data_counter[7]_net_1\, B => 
        \data_counter[8]_net_1\, Y => m27_m6_0_a2_4_2);
    
    \grant_counter_RNO[29]\ : XA1
      port map(A => \grant_counter[29]_net_1\, B => N_72, C => 
        N_202, Y => N_139);
    
    \DMAIn.Address[3]\ : DFN1E1C0
      port map(D => N_19, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[3]\);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_11 : NOR3C
      port map(A => \data_counter[27]_net_1\, B => 
        \data_counter[26]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_7_0, Y => 
        ADD_32x32_fast_I129_un1_Y_11_0);
    
    \state[1]\ : DFN1C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[1]_net_1\);
    
    un1_hresetn_inv_2_m30 : AX1C
      port map(A => \grant_counter[0]_net_1\, B => 
        un1_hresetn_inv_i_0, C => \grant_counter[1]_net_1\, Y => 
        N_31_0_i_0);
    
    \grant_counter_RNISQSF2[14]\ : OR3C
      port map(A => \state_ns_i_a2_0_i_o2_25[3]\, B => 
        \state_ns_i_a2_0_i_o2_24[3]\, C => 
        \state_ns_i_a2_0_i_o2_29[3]\, Y => N_246);
    
    \DMAIn.Burst\ : DFN1P0
      port map(D => N_194_i_0, CLK => HCLK_c, PRE => HRESETn_c, Q
         => Burst);
    
    un1_hresetn_inv_2_m18 : NOR3C
      port map(A => \grant_counter[2]_net_1\, B => N_17_0, C => 
        \grant_counter[3]_net_1\, Y => N_19_0);
    
    un1_hresetn_inv_2_m58 : AX1E
      port map(A => \grant_counter[21]_net_1\, B => N_56, C => 
        \grant_counter[22]_net_1\, Y => \un1_hresetn_inv_2_i[9]\);
    
    \data_counter_RNO[9]\ : XA1B
      port map(A => \data_counter[9]_net_1\, B => N_24_0_0, C => 
        N_198_0, Y => \data_counter_8[9]\);
    
    \DMAIn.Address_RNIK4FJ[17]\ : MX2
      port map(A => \Address[17]\, B => data_address(17), S => 
        time_select, Y => N_964);
    
    \data_counter_RNO[26]\ : XA1B
      port map(A => \data_counter[26]_net_1\, B => N_66, C => 
        N_198, Y => \data_counter_8[26]\);
    
    un1_hresetn_inv_2_m22 : NOR2B
      port map(A => N_22_0, B => \grant_counter[7]_net_1\, Y => 
        N_23_0);
    
    \state_RNO[3]\ : AO1C
      port map(A => N_241, B => N_235, C => \N_200\, Y => 
        \state_RNO[3]_net_1\);
    
    \state_RNO[0]\ : AO1D
      port map(A => N_241, B => N_235, C => 
        \state_RNO_0[0]_net_1\, Y => \state_RNO[0]_net_1\);
    
    \grant_counter[14]\ : DFN1
      port map(D => N_109, CLK => HCLK_c, Q => 
        \grant_counter[14]_net_1\);
    
    \grant_counter_RNICJK1[22]\ : NOR2B
      port map(A => \state_ns_i_a2_0_i_o2_22[3]\, B => 
        \state_ns_i_a2_0_i_o2_23[3]\, Y => 
        \state_ns_i_a2_0_i_o2_27[3]\);
    
    \DMAIn.Address[4]\ : DFN1E1C0
      port map(D => N_21, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[4]\);
    
    \grant_counter[2]\ : DFN1
      port map(D => \grant_counter_RNO[2]_net_1\, CLK => HCLK_c, 
        Q => \grant_counter[2]_net_1\);
    
    \data_counter_RNIB4B41[0]\ : MX2A
      port map(A => \state[5]_net_1\, B => 
        \data_counter[0]_net_1\, S => N_243, Y => N_508);
    
    \data_counter[26]\ : DFN1C0
      port map(D => \data_counter_8[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[26]_net_1\);
    
    \data_counter[23]\ : DFN1C0
      port map(D => \data_counter_8[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[23]_net_1\);
    
    \DMAIn.Address_RNIEIRJ[24]\ : MX2
      port map(A => \Address[24]\, B => data_address(24), S => 
        time_select_0, Y => N_971);
    
    \DMAIn.Address[25]\ : DFN1E1C0
      port map(D => N_69, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[25]\);
    
    un1_state_4_m45 : NOR3C
      port map(A => \data_counter[14]_net_1\, B => N623_0, C => 
        \data_counter[15]_net_1\, Y => N_46);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_8 : NOR3C
      port map(A => \data_counter[15]_net_1\, B => 
        \data_counter[14]_net_1\, C => 
        ADD_32x32_fast_I129_un1_Y_1_0, Y => 
        ADD_32x32_fast_I129_un1_Y_8_0);
    
    \grant_counter_RNO[19]\ : XA1
      port map(A => \grant_counter[19]_net_1\, B => N_52, C => 
        N_202, Y => N_119);
    
    \DMAIn.Address_RNO[2]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(2), Y
         => N_17);
    
    \data_counter_RNO[17]\ : XA1B
      port map(A => \data_counter[17]_net_1\, B => N_48_0, C => 
        N_198_0, Y => \data_counter_8[17]\);
    
    un1_state_4_m24 : NOR2B
      port map(A => N_24_0_0, B => \data_counter[9]_net_1\, Y => 
        N_25_0_0);
    
    \data_counter_RNO[25]\ : XA1B
      port map(A => \data_counter[25]_net_1\, B => N_64_0, C => 
        N_198, Y => \data_counter_8[25]\);
    
    \data_counter[21]\ : DFN1C0
      port map(D => \data_counter_8[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[21]_net_1\);
    
    \DMAIn.Address_RNO[4]\ : NOR2B
      port map(A => \state_0[5]_net_1\, B => data_address(4), Y
         => N_21);
    
    \grant_counter_RNO[7]\ : XA1
      port map(A => \grant_counter[7]_net_1\, B => N_22_0, C => 
        N_202_0, Y => N_95);
    
    \data_counter_RNI6F78[2]\ : NOR3C
      port map(A => \data_counter[2]_net_1\, B => 
        \data_counter[1]_net_1\, C => un1_state_5_i_o2_15, Y => 
        un1_state_5_i_o2_23);
    
    \DMAIn.Lock\ : DFN1E1C0
      port map(D => data_send, CLK => HCLK_c, CLR => HRESETn_c, E
         => \state[5]_net_1\, Q => Lock);
    
    \data_counter_RNO_3[0]\ : NOR2A
      port map(A => \state[0]_net_1\, B => 
        \data_counter[0]_net_1\, Y => N_337);
    
    \state_RNIQIK31_0[4]\ : OR2A
      port map(A => HRESETn_c, B => \N_200\, Y => N_202_0);
    
    \grant_counter[3]\ : DFN1
      port map(D => \grant_counter_RNO[3]_net_1\, CLK => HCLK_c, 
        Q => \grant_counter[3]_net_1\);
    
    \data_counter_RNIJUOF[10]\ : NOR2
      port map(A => \data_counter[10]_net_1\, B => 
        \data_counter[11]_net_1\, Y => un1_state_5_i_o2_5);
    
    \grant_counter[13]\ : DFN1
      port map(D => N_107, CLK => HCLK_c, Q => 
        \grant_counter[13]_net_1\);
    
    \grant_counter_RNIQOP[10]\ : NOR2B
      port map(A => \state_ns_i_a2_0_i_o2_6[3]\, B => 
        \state_ns_i_a2_0_i_o2_7[3]\, Y => 
        \state_ns_i_a2_0_i_o2_19[3]\);
    
    \grant_counter[27]\ : DFN1
      port map(D => N_135, CLK => HCLK_c, Q => 
        \grant_counter[27]_net_1\);
    
    \state_RNI1FH3[5]\ : NOR2B
      port map(A => \state[5]_net_1\, B => data_send, Y => 
        Request_5);
    
    \DMAIn.Address_RNIF4FJ[16]\ : MX2
      port map(A => \Address[16]\, B => data_address(16), S => 
        time_select, Y => N_963);
    
    \DMAIn.Address_RNIA4FJ[15]\ : MX2
      port map(A => \Address[15]\, B => data_address(15), S => 
        time_select, Y => N_962);
    
    un1_state_4_m15 : AOI1B
      port map(A => N_510, B => N_509, C => 
        \data_counter[0]_net_1\, Y => N_16_0);
    
    un1_hresetn_inv_2_m54 : AX1E
      port map(A => \grant_counter[19]_net_1\, B => N_52, C => 
        \grant_counter[20]_net_1\, Y => \un1_hresetn_inv_2_i[11]\);
    
    \grant_counter_RNIAQJD1[31]\ : NOR3C
      port map(A => \state_ns_i_a2_0_i_o2_3[3]\, B => 
        \state_ns_i_a2_0_i_o2_2[3]\, C => 
        \state_ns_i_a2_0_i_o2_16[3]\, Y => 
        \state_ns_i_a2_0_i_o2_24[3]\);
    
    \grant_counter[28]\ : DFN1
      port map(D => N_137, CLK => HCLK_c, Q => 
        \grant_counter[28]_net_1\);
    
    un1_state_4_ADD_32x32_fast_I174_Y_0 : XNOR2
      port map(A => N623_0, B => \data_counter[14]_net_1\, Y => 
        \un1_state_4_i[17]\);
    
    un1_hresetn_inv_2_m46 : AX1E
      port map(A => \grant_counter[15]_net_1\, B => N_44, C => 
        \grant_counter[16]_net_1\, Y => \un1_hresetn_inv_2_i[15]\);
    
    \grant_counter_RNIE9Q[22]\ : NOR3A
      port map(A => \state_ns_i_a2_0_i_o2_13[3]\, B => 
        \grant_counter[23]_net_1\, C => \grant_counter[22]_net_1\, 
        Y => \state_ns_i_a2_0_i_o2_22[3]\);
    
    \DMAIn.Address[26]\ : DFN1E1C0
      port map(D => N_71, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[26]\);
    
    \DMAIn.Address_RNIJ3361[6]\ : MX2
      port map(A => \Address[6]\, B => data_address(6), S => 
        time_select, Y => N_953);
    
    \data_counter_RNO[0]\ : NOR3
      port map(A => \data_counter_8_i_0[0]\, B => N_339, C => 
        N_336, Y => N_186);
    
    \state_RNIQ0SJ1[3]\ : NOR3B
      port map(A => HRESETn_c, B => Grant, C => N_241, Y => 
        un1_hresetn_inv_i_0);
    
    \state_RNIJBG8[0]\ : OR2B
      port map(A => \state[0]_net_1\, B => Ready, Y => N_346);
    
    \DMAIn.Address_RNIQHRJ[20]\ : MX2
      port map(A => \Address[20]\, B => data_address(20), S => 
        time_select_0, Y => N_967);
    
    \grant_counter_RNO[0]\ : AO1C
      port map(A => N_246, B => un1_hresetn_inv_i_0, C => 
        \grant_counter_0_0_0[0]\, Y => 
        \grant_counter_RNO[0]_net_1\);
    
    \data_counter[6]\ : DFN1C0
      port map(D => \data_counter_8[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[6]_net_1\);
    
    \data_counter[15]\ : DFN1C0
      port map(D => \data_counter_8[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[15]_net_1\);
    
    un1_state_4_ADD_32x32_fast_I129_un1_Y_3 : NOR2B
      port map(A => \data_counter[20]_net_1\, B => 
        \data_counter[21]_net_1\, Y => 
        ADD_32x32_fast_I129_un1_Y_3_0);
    
    un1_state_4_m47 : NOR2B
      port map(A => N_46, B => \data_counter[16]_net_1\, Y => 
        N_48_0);
    
    \data_counter_RNIDSMI6[22]\ : OR2B
      port map(A => un1_state_5_i_o2_30, B => un1_state_5_i_o2_29, 
        Y => N_235);
    
    un1_hresetn_inv_2_m63 : NOR3C
      port map(A => \grant_counter[23]_net_1\, B => N_60, C => 
        \grant_counter[24]_net_1\, Y => N_64);
    
    \data_counter_RNO[19]\ : XA1B
      port map(A => \data_counter[19]_net_1\, B => N_52_0, C => 
        N_198_0, Y => \data_counter_8[19]\);
    
    \grant_counter_RNO[8]\ : XA1
      port map(A => \grant_counter[8]_net_1\, B => N_23_0, C => 
        N_202_0, Y => N_97);
    
    \data_counter[20]\ : DFN1C0
      port map(D => \data_counter_8[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[20]_net_1\);
    
    un1_state_4_m28_m6 : NOR3B
      port map(A => m28_m6_5, B => m27_m6_0_a2_4, C => N_243, Y
         => N623_0);
    
    un1_hresetn_inv_2_ADD_32x32_fast_I129_un1_Y_13 : NOR3C
      port map(A => ADD_32x32_fast_I129_un1_Y_5, B => 
        ADD_32x32_fast_I129_un1_Y_4, C => 
        ADD_32x32_fast_I129_un1_Y_11, Y => 
        ADD_32x32_fast_I129_un1_Y_13);
    
    \data_counter[22]\ : DFN1C0
      port map(D => \data_counter_8[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_counter[22]_net_1\);
    
    \data_counter_RNIQDKV[15]\ : NOR3A
      port map(A => un1_state_5_i_o2_7, B => 
        \data_counter[15]_net_1\, C => \data_counter[14]_net_1\, 
        Y => un1_state_5_i_o2_19);
    
    \state_RNIU9K11[4]\ : AO1C
      port map(A => Grant, B => \state[4]_net_1\, C => 
        un1_state_2_i_o2_0, Y => N_243);
    
    \grant_counter_RNIAPP[14]\ : NOR3A
      port map(A => \state_ns_i_a2_0_i_o2_9[3]\, B => 
        \grant_counter[15]_net_1\, C => \grant_counter[14]_net_1\, 
        Y => \state_ns_i_a2_0_i_o2_20[3]\);
    
    \DMAIn.Address[27]\ : DFN1E1C0
      port map(D => N_73, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_154, Q => \Address[27]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\ is

    port( nb_burst_available  : in    std_logic_vector(10 downto 0);
          status_full_err     : out   std_logic_vector(1 to 1);
          status_full         : out   std_logic_vector(1 to 1);
          sel_data            : in    std_logic_vector(1 to 1);
          sel_data_0          : in    std_logic_vector(1 to 1);
          update_and_sel_5    : in    std_logic_vector(3 downto 2);
          addr_data_f1        : in    std_logic_vector(31 downto 0);
          status_full_ack     : in    std_logic_vector(1 to 1);
          addr_data_vector_94 : in    std_logic;
          addr_data_vector_91 : in    std_logic;
          addr_data_vector_89 : in    std_logic;
          addr_data_vector_87 : in    std_logic;
          addr_data_vector_86 : in    std_logic;
          addr_data_vector_85 : in    std_logic;
          addr_data_vector_84 : in    std_logic;
          addr_data_vector_83 : in    std_logic;
          addr_data_vector_67 : in    std_logic;
          addr_data_vector_66 : in    std_logic;
          addr_data_vector_65 : in    std_logic;
          addr_data_vector_64 : in    std_logic;
          addr_data_vector_75 : in    std_logic;
          addr_data_vector_73 : in    std_logic;
          addr_data_vector_81 : in    std_logic;
          addr_data_vector_79 : in    std_logic;
          addr_data_vector_77 : in    std_logic;
          addr_data_vector_24 : out   std_logic;
          addr_data_vector_31 : out   std_logic;
          addr_data_vector_16 : out   std_logic;
          addr_data_vector_14 : out   std_logic;
          addr_data_vector_18 : out   std_logic;
          addr_data_vector_26 : out   std_logic;
          addr_data_vector_29 : out   std_logic;
          addr_data_vector_28 : out   std_logic;
          addr_data_vector_5  : out   std_logic;
          addr_data_vector_4  : out   std_logic;
          addr_data_vector_6  : out   std_logic;
          addr_data_vector_12 : out   std_logic;
          addr_data_vector_10 : out   std_logic;
          addr_data_vector_7  : out   std_logic;
          addr_data_vector_8  : out   std_logic;
          N_913               : out   std_logic;
          N_910               : out   std_logic;
          N_908               : out   std_logic;
          N_906               : out   std_logic;
          N_905               : out   std_logic;
          N_904               : out   std_logic;
          N_903               : out   std_logic;
          N_902               : out   std_logic;
          N_1300              : out   std_logic;
          N_1299              : out   std_logic;
          N_1298              : out   std_logic;
          N_1297              : out   std_logic;
          N_1294              : out   std_logic;
          N_1292              : out   std_logic;
          N_1286              : out   std_logic;
          N_1284              : out   std_logic;
          N_1282              : out   std_logic;
          HRESETn_c           : in    std_logic;
          HCLK_c              : in    std_logic
        );

end 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\ is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \state_0[0]_net_1\, N_118, N_38, \nb_send[1]_net_1\, 
        \nb_send[0]_net_1\, N_30, \nb_send[3]_net_1\, 
        \DWACT_FINC_E[0]\, N_7, \nb_send[8]_net_1\, 
        \DWACT_FINC_E[4]\, m40_m6_0_a2_6, m40_m6_0_a2_1, 
        m40_m6_0_a2_0, m40_m6_0_a2_5, m40_m6_0_a2_3, 
        \addr_data_vector[41]\, \addr_data_vector[54]\, 
        \addr_data_vector[55]\, \addr_data_vector[43]\, 
        m20_m7_i_4, address_0_sqmuxa, m20_m7_i_3, m20_m7_i_0, 
        \addr_data_vector[42]\, m20_m7_i_1, 
        \addr_data_vector[40]\, \addr_data_vector[39]\, 
        m20_m3_e_0, \un1_state_12_3_0[4]\, \update_r_i[0]\, 
        \update_r[1]_net_1\, address_0_sqmuxa_0, \state[3]_net_1\, 
        un3_update_r, un1_state_5_i_0, \state[4]_net_1\, 
        \state_ns_i_0[3]\, N_131, address_7_31_m6_e_3, 
        \addr_data_vector[57]\, \addr_data_vector[62]\, 
        address_7_31_m6_e_1, address_7_31_m6_e_2, 
        \addr_data_vector[59]\, m36_m6_0_a2_4_6, 
        \addr_data_vector[51]\, m36_m6_0_a2_4_4, m36_m6_0_a2_4_5, 
        \addr_data_vector[47]\, m36_m6_0_a2_4_2, 
        \addr_data_vector[45]\, \addr_data_vector[53]\, 
        \addr_data_vector[52]\, \addr_data_vector[49]\, 
        \un1_address[6]\, \addr_data_vector[38]\, N_5_0, N_116, 
        N_129, \state[1]_net_1\, \state_ns[0]\, N_125, N_124, 
        \un1_state_12_2[4]\, N_110, \state[2]_net_1\, state7, 
        m36_m6_0_a2_4_i, \address_RNO_2[31]_net_1\, N_41, N_13_0, 
        m20_m3_e, N_69, m20_N_17_i_0, m20_m7_i_o5, 
        \address_7[31]\, \address_RNO_0[31]_net_1\, 
        \address_RNO_1[31]_net_1\, \addr_data_vector[63]\, N_37_0, 
        \addr_data_vector[44]\, N_2, \addr_data_vector[34]\, 
        N_15_0_i_0, N_16_0, N_17_0_i_0, N_18_0, N_20_0_i_0, 
        N_22_0_i_0, N_24_0, N_26_0_i_0, \addr_data_vector[46]\, 
        N_27_0, N_28_0_i_0, \addr_data_vector[48]\, N_30_0_i_0, 
        N_31_0, \un1_address[19]\, \addr_data_vector[50]\, N_34_0, 
        \un1_address[20]\, \un1_address[23]\, N_40_i_0, N_43, 
        \addr_data_vector[56]\, N_45, \addr_data_vector[58]\, 
        N_46, \addr_data_vector[60]\, N_50_i_0, 
        \addr_data_vector[35]\, N_51_i_0, \addr_data_vector[36]\, 
        N_52_i_0, \addr_data_vector[37]\, N_1_i_0, N_54_0_i_0, 
        N_55_0_i_0, \un1_address[18]\, \un1_address[21]\, 
        \un1_address[22]\, \un1_address[24]\, \un1_address[25]\, 
        \un1_address[26]\, \un1_address[27]\, \un1_address[28]\, 
        \un1_address[29]\, \addr_data_vector[61]\, 
        \un1_address[30]\, \address_7[2]\, \address_7[3]\, 
        \address_7[4]\, \address_7[5]\, \address_7[6]\, 
        \address_7[7]\, \address_7[8]\, \address_7[9]\, 
        \address_7[10]\, \address_7[11]\, \address_7[12]\, 
        \address_7[13]\, \address_7[15]\, \address_7[16]\, 
        \address_7[17]\, \state[0]_net_1\, \address_7[18]\, 
        \address_7[19]\, \address_7[20]\, \address_7[21]\, 
        \address_7[22]\, \address_7[23]\, \address_7[24]\, 
        \address_7[25]\, \address_7[26]\, \address_7[27]\, 
        \address_7[28]\, \address_7[29]\, \address_7[30]\, 
        N_56_0_i_0, un1_state_9, \nb_send_5[0]\, \nb_send_5[1]\, 
        \un2_nb_send_next[1]\, \nb_send_5[2]\, 
        \un2_nb_send_next[2]\, \nb_send_5[3]\, 
        \un2_nb_send_next[3]\, \nb_send_5[4]\, 
        \un2_nb_send_next[4]\, \nb_send_5[5]\, 
        \un2_nb_send_next[5]\, \nb_send_5[6]\, 
        \un2_nb_send_next[6]\, \nb_send_5[7]\, 
        \un2_nb_send_next[7]\, \nb_send_5[8]\, 
        \un2_nb_send_next[8]\, \nb_send_5[9]\, 
        \un2_nb_send_next[9]\, \nb_send_5[10]\, 
        \un2_nb_send_next[10]\, N_127, N_113, \state_ns[2]\, 
        un1_state_11, \address_7[14]\, \addr_data_vector[32]\, 
        \addr_data_vector[33]\, \nb_send[2]_net_1\, 
        \nb_send[4]_net_1\, \nb_send[5]_net_1\, 
        \nb_send[6]_net_1\, \nb_send[7]_net_1\, 
        \nb_send[9]_net_1\, \nb_send[10]_net_1\, N_4, 
        \DWACT_FINC_E[2]\, \DWACT_FINC_E[3]\, N_12, N_17, N_22, 
        \DWACT_FINC_E[1]\, N_27, N_35, \DWACT_COMP0_E[1]\, 
        \DWACT_COMP0_E[2]\, \DWACT_COMP0_E[0]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, \ACT_LT4_E[3]\, 
        \ACT_LT4_E[6]\, \ACT_LT4_E[10]\, \ACT_LT4_E[7]\, 
        \ACT_LT4_E[8]\, \ACT_LT4_E[5]\, \ACT_LT4_E[4]\, 
        \ACT_LT4_E[0]\, \ACT_LT4_E[1]\, \ACT_LT4_E[2]\, 
        \ACT_LT2_E[0]\, \ACT_LT2_E[1]\, \ACT_LT2_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, N_37, 
        N_36, N_35_0, N_32, N_34, N_33, N_31, N_28, N_29, N_30_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, 
        \DWACT_BL_EQUAL_0_E[4]\, \DWACT_BL_EQUAL_0_E[3]\, 
        \DWACT_BL_EQUAL_0_E_0[0]\, \DWACT_BL_EQUAL_0_E_0[1]\, 
        \DWACT_BL_EQUAL_0_E[2]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    addr_data_vector_24 <= \addr_data_vector[56]\;
    addr_data_vector_31 <= \addr_data_vector[63]\;
    addr_data_vector_16 <= \addr_data_vector[48]\;
    addr_data_vector_14 <= \addr_data_vector[46]\;
    addr_data_vector_18 <= \addr_data_vector[50]\;
    addr_data_vector_26 <= \addr_data_vector[58]\;
    addr_data_vector_29 <= \addr_data_vector[61]\;
    addr_data_vector_28 <= \addr_data_vector[60]\;
    addr_data_vector_5 <= \addr_data_vector[37]\;
    addr_data_vector_4 <= \addr_data_vector[36]\;
    addr_data_vector_6 <= \addr_data_vector[38]\;
    addr_data_vector_12 <= \addr_data_vector[44]\;
    addr_data_vector_10 <= \addr_data_vector[42]\;
    addr_data_vector_7 <= \addr_data_vector[39]\;
    addr_data_vector_8 <= \addr_data_vector[40]\;

    \address[16]\ : DFN1C0
      port map(D => \address_7[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[48]\);
    
    \address[10]\ : DFN1C0
      port map(D => \address_7[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[42]\);
    
    \state[0]\ : DFN1C0
      port map(D => N_118, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[0]_net_1\);
    
    \address[30]\ : DFN1C0
      port map(D => \address_7[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[62]\);
    
    un1_address_m20_m7_i_0 : NOR2B
      port map(A => \addr_data_vector[43]\, B => 
        \addr_data_vector[39]\, Y => m20_m7_i_0);
    
    un1_address_m45 : NOR2A
      port map(A => \addr_data_vector[60]\, B => N_45, Y => N_46);
    
    \address_RNO[26]\ : MX2
      port map(A => \un1_address[26]\, B => addr_data_f1(26), S
         => \state[0]_net_1\, Y => \address_7[26]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_25\ : AO1C
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_31, Y => N_36);
    
    un1_address_m61 : XNOR2
      port map(A => N_43, B => \addr_data_vector[58]\, Y => 
        \un1_address[26]\);
    
    \address[26]\ : DFN1C0
      port map(D => \address_7[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[58]\);
    
    \address[20]\ : DFN1C0
      port map(D => \address_7[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[52]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_42\ : AO1C
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => \un2_nb_send_next[5]\, Y => 
        \ACT_LT2_E[1]\);
    
    \state_RNO_0[2]\ : NOR3B
      port map(A => N_129, B => \state[2]_net_1\, C => 
        status_full_ack(1), Y => N_127);
    
    \state_RNI3CSP8[3]\ : OR2B
      port map(A => \state[3]_net_1\, B => state7, Y => 
        \un1_state_12_2[4]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_57\ : NOR2A
      port map(A => \ACT_LT4_E[4]\, B => \ACT_LT4_E[5]\, Y => 
        \ACT_LT4_E[6]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_36\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[1]\, B => 
        \DWACT_BL_EQUAL_0_E[0]\, Y => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\);
    
    un1_address_m51 : AX1C
      port map(A => \addr_data_vector[36]\, B => N_69, C => 
        \addr_data_vector[37]\, Y => N_52_i_0);
    
    \address[12]\ : DFN1C0
      port map(D => \address_7[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[44]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_22\ : OA1A
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), C => N_29, Y => N_33);
    
    \address_RNO[29]\ : MX2
      port map(A => \un1_address[29]\, B => addr_data_f1(29), S
         => \state[0]_net_1\, Y => \address_7[29]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_8\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, B => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, Y => 
        \DWACT_COMP0_E[1]\);
    
    un1_address_m36_m6_0_a2_4_4 : NOR3C
      port map(A => \addr_data_vector[45]\, B => 
        \addr_data_vector[53]\, C => \addr_data_vector[52]\, Y
         => m36_m6_0_a2_4_4);
    
    un1_address_m36_m6_0_a2_4 : OR2B
      port map(A => m36_m6_0_a2_4_6, B => m36_m6_0_a2_4_5, Y => 
        m36_m6_0_a2_4_i);
    
    un1_address_m19 : AX1C
      port map(A => \addr_data_vector[42]\, B => N_18_0, C => 
        \addr_data_vector[43]\, Y => N_20_0_i_0);
    
    \address_RNI68OA[9]\ : MX2C
      port map(A => \addr_data_vector[41]\, B => 
        addr_data_vector_73, S => sel_data_0(1), Y => N_1292);
    
    \address[22]\ : DFN1C0
      port map(D => \address_7[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[54]\);
    
    \address_RNO[23]\ : MX2
      port map(A => \un1_address[23]\, B => addr_data_f1(23), S
         => \state[0]_net_1\, Y => \address_7[23]\);
    
    \address[2]\ : DFN1C0
      port map(D => \address_7[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[34]\);
    
    un2_nb_send_next_I_13 : XOR2
      port map(A => N_35, B => \nb_send[3]_net_1\, Y => 
        \un2_nb_send_next[3]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_54\ : AOI1A
      port map(A => \ACT_LT4_E[0]\, B => \ACT_LT4_E[1]\, C => 
        \ACT_LT4_E[2]\, Y => \ACT_LT4_E[3]\);
    
    \address_RNO[24]\ : MX2
      port map(A => \un1_address[24]\, B => addr_data_f1(24), S
         => \state[0]_net_1\, Y => \address_7[24]\);
    
    \address_RNO[10]\ : MX2
      port map(A => N_54_0_i_0, B => addr_data_f1(10), S => 
        \state_0[0]_net_1\, Y => \address_7[10]\);
    
    \status_full_err\ : DFN1E0C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_110, Q => status_full_err(1));
    
    un2_nb_send_next_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \nb_send[8]_net_1\, C
         => \nb_send[9]_net_1\, Y => N_4);
    
    \nb_send_RNO[1]\ : NOR2B
      port map(A => \un2_nb_send_next[1]\, B => state7, Y => 
        \nb_send_5[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_51\ : NOR2B
      port map(A => \nb_send[0]_net_1\, B => 
        nb_burst_available(0), Y => \ACT_LT4_E[0]\);
    
    un2_nb_send_next_I_31 : XOR2
      port map(A => N_22, B => \nb_send[6]_net_1\, Y => 
        \un2_nb_send_next[6]\);
    
    \nb_send[9]\ : DFN1E0C0
      port map(D => \nb_send_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[9]_net_1\);
    
    \address_RNO[9]\ : MX2
      port map(A => N_17_0_i_0, B => addr_data_f1(9), S => 
        \state_0[0]_net_1\, Y => \address_7[9]\);
    
    \address[5]\ : DFN1C0
      port map(D => \address_7[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[37]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_5\ : XNOR2
      port map(A => \un2_nb_send_next[7]\, B => 
        nb_burst_available(7), Y => \DWACT_BL_EQUAL_0_E_0[1]\);
    
    \address[15]\ : DFN1C0
      port map(D => \address_7[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[47]\);
    
    \address[13]\ : DFN1C0
      port map(D => \address_7[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[45]\);
    
    \state[4]\ : DFN1P0
      port map(D => \state_ns[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[4]_net_1\);
    
    \nb_send_RNO[9]\ : NOR2B
      port map(A => \un2_nb_send_next[9]\, B => state7, Y => 
        \nb_send_5[9]\);
    
    \address[19]\ : DFN1C0
      port map(D => \address_7[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[51]\);
    
    \address[25]\ : DFN1C0
      port map(D => \address_7[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[57]\);
    
    un2_nb_send_next_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => \nb_send[5]_net_1\, Y => N_22);
    
    \address[23]\ : DFN1C0
      port map(D => \address_7[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[55]\);
    
    un1_address_m14 : AX1
      port map(A => N_13_0, B => \addr_data_vector[39]\, C => 
        \addr_data_vector[40]\, Y => N_15_0_i_0);
    
    un1_address_m29 : AX1C
      port map(A => \addr_data_vector[48]\, B => N_27_0, C => 
        \addr_data_vector[49]\, Y => N_30_0_i_0);
    
    un2_nb_send_next_I_12 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => N_35);
    
    \FSM_SELECT_ADDRESS.state7_0_I_19\ : NOR2A
      port map(A => nb_burst_available(6), B => 
        \un2_nb_send_next[6]\, Y => N_30_0);
    
    un1_address_m36_m6_0_a2 : NOR3B
      port map(A => \addr_data_vector[44]\, B => m20_N_17_i_0, C
         => m36_m6_0_a2_4_i, Y => N_37_0);
    
    \address_RNO_2[31]\ : NOR3B
      port map(A => address_7_31_m6_e_3, B => address_7_31_m6_e_2, 
        C => \state_0[0]_net_1\, Y => \address_RNO_2[31]_net_1\);
    
    \address[29]\ : DFN1C0
      port map(D => \address_7[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[61]\);
    
    \address[18]\ : DFN1C0
      port map(D => \address_7[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[50]\);
    
    \nb_send_RNO[6]\ : NOR2B
      port map(A => \un2_nb_send_next[6]\, B => state7, Y => 
        \nb_send_5[6]\);
    
    \address_RNO[21]\ : MX2
      port map(A => \un1_address[21]\, B => addr_data_f1(21), S
         => \state[0]_net_1\, Y => \address_7[21]\);
    
    \address_RNO[16]\ : MX2
      port map(A => N_28_0_i_0, B => addr_data_f1(16), S => 
        \state_0[0]_net_1\, Y => \address_7[16]\);
    
    un2_nb_send_next_I_51 : NOR2B
      port map(A => \nb_send[8]_net_1\, B => \DWACT_FINC_E[4]\, Y
         => N_7);
    
    \address[0]\ : DFN1E1C0
      port map(D => addr_data_f1(0), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        \addr_data_vector[32]\);
    
    status_full_err_RNO_0 : OR2
      port map(A => \state[4]_net_1\, B => \state[3]_net_1\, Y
         => un1_state_5_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_address_m36_m6_0_a2_4_2 : NOR2B
      port map(A => \addr_data_vector[48]\, B => 
        \addr_data_vector[49]\, Y => m36_m6_0_a2_4_2);
    
    \address_RNO[27]\ : MX2
      port map(A => \un1_address[27]\, B => addr_data_f1(27), S
         => \state[0]_net_1\, Y => \address_7[27]\);
    
    \address[4]\ : DFN1C0
      port map(D => \address_7[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[36]\);
    
    \address[28]\ : DFN1C0
      port map(D => \address_7[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[60]\);
    
    un1_address_m1 : NOR3A
      port map(A => \addr_data_vector[34]\, B => 
        \un1_state_12_2[4]\, C => \un1_state_12_3_0[4]\, Y => N_2);
    
    \FSM_SELECT_ADDRESS.state7_0_I_7\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[4]\, B => 
        \DWACT_BL_EQUAL_0_E[3]\, Y => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\);
    
    un1_address_m17 : NOR2A
      port map(A => \addr_data_vector[41]\, B => N_16_0, Y => 
        N_18_0);
    
    \nb_send_RNO[2]\ : NOR2B
      port map(A => \un2_nb_send_next[2]\, B => state7, Y => 
        \nb_send_5[2]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \state_RNO_0[4]\ : OR3B
      port map(A => N_131, B => N_129, C => \state[3]_net_1\, Y
         => N_125);
    
    \address_RNO_1[31]\ : AX1E
      port map(A => \addr_data_vector[56]\, B => N_41, C => 
        \addr_data_vector[63]\, Y => \address_RNO_1[31]_net_1\);
    
    un1_address_m20_m7_i_4 : OA1A
      port map(A => address_0_sqmuxa, B => \addr_data_vector[38]\, 
        C => m20_m7_i_3, Y => m20_m7_i_4);
    
    \FSM_SELECT_ADDRESS.state7_0_I_58\ : NOR2A
      port map(A => \un2_nb_send_next[2]\, B => 
        nb_burst_available(2), Y => \ACT_LT4_E[7]\);
    
    \nb_send_RNO[7]\ : NOR2B
      port map(A => \un2_nb_send_next[7]\, B => state7, Y => 
        \nb_send_5[7]\);
    
    un2_nb_send_next_I_24 : XOR2
      port map(A => N_27, B => \nb_send[5]_net_1\, Y => 
        \un2_nb_send_next[5]\);
    
    un2_nb_send_next_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \nb_send[3]_net_1\, C
         => \nb_send[4]_net_1\, Y => N_27);
    
    un1_address_ADD_32x32_fast_I164_Y_0 : XOR3
      port map(A => address_0_sqmuxa, B => \addr_data_vector[38]\, 
        C => N_5_0, Y => \un1_address[6]\);
    
    \address_RNO[19]\ : MX2
      port map(A => \un1_address[19]\, B => addr_data_f1(19), S
         => \state[0]_net_1\, Y => \address_7[19]\);
    
    \nb_send[7]\ : DFN1E0C0
      port map(D => \nb_send_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[7]_net_1\);
    
    un1_address_m40_m6_0_a2_5 : NOR3C
      port map(A => \addr_data_vector[40]\, B => 
        \addr_data_vector[39]\, C => m40_m6_0_a2_3, Y => 
        m40_m6_0_a2_5);
    
    \address_RNO[13]\ : MX2
      port map(A => N_55_0_i_0, B => addr_data_f1(13), S => 
        \state_0[0]_net_1\, Y => \address_7[13]\);
    
    \address_RNIFA45[30]\ : MX2C
      port map(A => \addr_data_vector[62]\, B => 
        addr_data_vector_94, S => sel_data(1), Y => N_913);
    
    \address[14]\ : DFN1C0
      port map(D => \address_7[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[46]\);
    
    \state_RNO[1]\ : OA1C
      port map(A => N_129, B => \state[1]_net_1\, C => 
        \state_ns_i_0[3]\, Y => N_116);
    
    \nb_send[0]\ : DFN1E0C0
      port map(D => \nb_send_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[0]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_53\ : AND2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[2]\);
    
    \address_RNIJ245[25]\ : MX2C
      port map(A => \addr_data_vector[57]\, B => 
        addr_data_vector_89, S => sel_data(1), Y => N_908);
    
    \nb_send[6]\ : DFN1E0C0
      port map(D => \nb_send_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[6]_net_1\);
    
    \nb_send[10]\ : DFN1E0C0
      port map(D => \nb_send_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[10]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_56\ : NOR2A
      port map(A => nb_burst_available(3), B => 
        \un2_nb_send_next[3]\, Y => \ACT_LT4_E[5]\);
    
    \address_RNO[14]\ : MX2
      port map(A => N_56_0_i_0, B => addr_data_f1(14), S => 
        \state[0]_net_1\, Y => \address_7[14]\);
    
    un1_address_m20_m3_e_0 : NOR2B
      port map(A => \addr_data_vector[36]\, B => 
        \addr_data_vector[37]\, Y => m20_m3_e_0);
    
    \nb_send_RNO[3]\ : NOR2B
      port map(A => \un2_nb_send_next[3]\, B => state7, Y => 
        \nb_send_5[3]\);
    
    \nb_send[2]\ : DFN1E0C0
      port map(D => \nb_send_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[2]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_27\ : OA1
      port map(A => N_37, B => N_36, C => N_35_0, Y => 
        \DWACT_COMP0_E[0]\);
    
    \address[24]\ : DFN1C0
      port map(D => \address_7[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[56]\);
    
    un1_address_m27 : XOR2
      port map(A => N_27_0, B => \addr_data_vector[48]\, Y => 
        N_28_0_i_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \address_RNO_0[31]\ : MX2C
      port map(A => \addr_data_vector[63]\, B => addr_data_f1(31), 
        S => \state_0[0]_net_1\, Y => \address_RNO_0[31]_net_1\);
    
    \address_RNILQ35[19]\ : MX2C
      port map(A => \addr_data_vector[51]\, B => 
        addr_data_vector_83, S => sel_data(1), Y => N_902);
    
    un1_address_m60 : AX1C
      port map(A => \addr_data_vector[56]\, B => N_41, C => 
        \addr_data_vector[57]\, Y => \un1_address[25]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_44\ : AND3A
      port map(A => \ACT_LT2_E[0]\, B => \ACT_LT2_E[1]\, C => 
        \ACT_LT2_E[2]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\);
    
    un1_address_m36_m6_0_a2_4_5 : NOR3C
      port map(A => \addr_data_vector[47]\, B => 
        \addr_data_vector[46]\, C => m36_m6_0_a2_4_2, Y => 
        m36_m6_0_a2_4_5);
    
    un1_address_m30 : NOR3C
      port map(A => \addr_data_vector[48]\, B => N_27_0, C => 
        \addr_data_vector[49]\, Y => N_31_0);
    
    \nb_send[4]\ : DFN1E0C0
      port map(D => \nb_send_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[4]_net_1\);
    
    un1_address_m16 : XNOR2
      port map(A => N_16_0, B => \addr_data_vector[41]\, Y => 
        N_17_0_i_0);
    
    un2_nb_send_next_I_45 : XOR2
      port map(A => N_12, B => \nb_send[8]_net_1\, Y => 
        \un2_nb_send_next[8]\);
    
    \nb_send_RNO[0]\ : NOR2A
      port map(A => state7, B => \nb_send[0]_net_1\, Y => 
        \nb_send_5[0]\);
    
    \nb_send_RNO[8]\ : NOR2B
      port map(A => \un2_nb_send_next[8]\, B => state7, Y => 
        \nb_send_5[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_41\ : AND2A
      port map(A => nb_burst_available(5), B => 
        \un2_nb_send_next[5]\, Y => \ACT_LT2_E[0]\);
    
    \state_RNO[4]\ : OR3C
      port map(A => N_125, B => N_124, C => \un1_state_12_2[4]\, 
        Y => \state_ns[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_4\ : XNOR2
      port map(A => \un2_nb_send_next[9]\, B => 
        nb_burst_available(9), Y => \DWACT_BL_EQUAL_0_E[3]\);
    
    \address[8]\ : DFN1C0
      port map(D => \address_7[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[40]\);
    
    un1_address_m50 : XOR2
      port map(A => N_69, B => \addr_data_vector[36]\, Y => 
        N_51_i_0);
    
    un1_address_m39 : AX1B
      port map(A => \un1_state_12_2[4]\, B => 
        \un1_state_12_3_0[4]\, C => \addr_data_vector[34]\, Y => 
        N_40_i_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_24\ : OR2A
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => N_35_0);
    
    \state_ns_i_a2[1]\ : NOR2A
      port map(A => update_and_sel_5(2), B => update_and_sel_5(3), 
        Y => N_129);
    
    \address_RNO[6]\ : MX2
      port map(A => \un1_address[6]\, B => addr_data_f1(6), S => 
        \state_0[0]_net_1\, Y => \address_7[6]\);
    
    \state_RNO[2]\ : AO1A
      port map(A => state7, B => \state[3]_net_1\, C => N_127, Y
         => \state_ns[2]\);
    
    \address_RNO[28]\ : MX2
      port map(A => \un1_address[28]\, B => addr_data_f1(28), S
         => \state[0]_net_1\, Y => \address_7[28]\);
    
    \address_RNO[11]\ : MX2
      port map(A => N_20_0_i_0, B => addr_data_f1(11), S => 
        \state_0[0]_net_1\, Y => \address_7[11]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_21\ : AO1C
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, C => N_30_0, Y => N_32);
    
    un1_address_m40_m6_0_a2_3 : NOR2B
      port map(A => \addr_data_vector[41]\, B => 
        \addr_data_vector[42]\, Y => m40_m6_0_a2_3);
    
    \FSM_SELECT_ADDRESS.state7_0_I_73\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => state7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_35\ : XNOR2
      port map(A => \un2_nb_send_next[5]\, B => 
        nb_burst_available(5), Y => \DWACT_BL_EQUAL_0_E[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_2\ : XNOR2
      port map(A => \un2_nb_send_next[6]\, B => 
        nb_burst_available(6), Y => \DWACT_BL_EQUAL_0_E_0[0]\);
    
    un1_address_m38 : AX1C
      port map(A => \addr_data_vector[54]\, B => N_37_0, C => 
        \addr_data_vector[55]\, Y => \un1_address[23]\);
    
    un1_address_m12 : AO13
      port map(A => N_5_0, B => address_0_sqmuxa, C => 
        \addr_data_vector[38]\, Y => N_13_0);
    
    un1_address_m59 : XOR2
      port map(A => N_41, B => \addr_data_vector[56]\, Y => 
        \un1_address[24]\);
    
    \address_RNIB245[21]\ : MX2C
      port map(A => \addr_data_vector[53]\, B => 
        addr_data_vector_85, S => sel_data(1), Y => N_904);
    
    \update_r[0]\ : DFN1P0
      port map(D => update_and_sel_5(2), CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \update_r_i[0]\);
    
    un2_nb_send_next_I_5 : XOR2
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        Y => \un2_nb_send_next[1]\);
    
    un1_address_m40_m6_0_a2_6 : NOR3C
      port map(A => m40_m6_0_a2_1, B => m40_m6_0_a2_0, C => 
        m40_m6_0_a2_5, Y => m40_m6_0_a2_6);
    
    \address_RNO[17]\ : MX2
      port map(A => N_30_0_i_0, B => addr_data_f1(17), S => 
        \state[0]_net_1\, Y => \address_7[17]\);
    
    \address_RNO[5]\ : MX2
      port map(A => N_52_i_0, B => addr_data_f1(5), S => 
        \state_0[0]_net_1\, Y => \address_7[5]\);
    
    un1_address_m15 : OR3B
      port map(A => \addr_data_vector[39]\, B => 
        \addr_data_vector[40]\, C => N_13_0, Y => N_16_0);
    
    un1_address_m58 : XOR2
      port map(A => N_37_0, B => \addr_data_vector[54]\, Y => 
        \un1_address[22]\);
    
    \state_RNI40SU8[3]\ : AO1B
      port map(A => un3_update_r, B => state7, C => 
        \state[3]_net_1\, Y => un1_state_9);
    
    un2_nb_send_next_I_56 : XOR2
      port map(A => N_4, B => \nb_send[10]_net_1\, Y => 
        \un2_nb_send_next[10]\);
    
    un1_address_m26 : NOR3C
      port map(A => \addr_data_vector[46]\, B => N_24_0, C => 
        \addr_data_vector[47]\, Y => N_27_0);
    
    un2_nb_send_next_I_41 : AND2
      port map(A => \nb_send[6]_net_1\, B => \nb_send[7]_net_1\, 
        Y => \DWACT_FINC_E[3]\);
    
    \address_RNO[3]\ : MX2
      port map(A => N_50_i_0, B => addr_data_f1(3), S => 
        \state_0[0]_net_1\, Y => \address_7[3]\);
    
    \address_RNO_4[31]\ : NOR2B
      port map(A => \addr_data_vector[60]\, B => 
        \addr_data_vector[61]\, Y => address_7_31_m6_e_2);
    
    \address[3]\ : DFN1C0
      port map(D => \address_7[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[35]\);
    
    un2_nb_send_next_I_34 : AND3
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        C => \nb_send[5]_net_1\, Y => \DWACT_FINC_E[2]\);
    
    un1_address_m64 : XOR2
      port map(A => N_46, B => \addr_data_vector[61]\, Y => 
        \un1_address[29]\);
    
    un1_address_m34 : XOR2
      port map(A => N_34_0, B => \addr_data_vector[52]\, Y => 
        \un1_address[20]\);
    
    \address_RNO[30]\ : MX2
      port map(A => \un1_address[30]\, B => addr_data_f1(30), S
         => \state[0]_net_1\, Y => \address_7[30]\);
    
    \address_RNI9245[20]\ : MX2C
      port map(A => \addr_data_vector[52]\, B => 
        addr_data_vector_84, S => sel_data(1), Y => N_903);
    
    \state_RNO_0[1]\ : OR2
      port map(A => status_full_ack(1), B => N_131, Y => 
        \state_ns_i_0[3]\);
    
    \state_RNITJCD[1]\ : NOR2
      port map(A => \state[2]_net_1\, B => \state[1]_net_1\, Y
         => N_131);
    
    \nb_send[3]\ : DFN1E0C0
      port map(D => \nb_send_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[3]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_20\ : OR2A
      port map(A => nb_burst_available(10), B => 
        \un2_nb_send_next[10]\, Y => N_31);
    
    un1_address_m54 : AX1C
      port map(A => \addr_data_vector[44]\, B => m20_N_17_i_0, C
         => \addr_data_vector[45]\, Y => N_55_0_i_0);
    
    \address[7]\ : DFN1C0
      port map(D => \address_7[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[39]\);
    
    un2_nb_send_next_I_38 : XOR2
      port map(A => N_17, B => \nb_send[7]_net_1\, Y => 
        \un2_nb_send_next[7]\);
    
    \nb_send[5]\ : DFN1E0C0
      port map(D => \nb_send_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[5]_net_1\);
    
    \nb_send_RNO[5]\ : NOR2B
      port map(A => \un2_nb_send_next[5]\, B => state7, Y => 
        \nb_send_5[5]\);
    
    un1_address_m25 : AX1C
      port map(A => \addr_data_vector[46]\, B => N_24_0, C => 
        \addr_data_vector[47]\, Y => N_26_0_i_0);
    
    \state[3]\ : DFN1C0
      port map(D => N_113, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[3]_net_1\);
    
    \address_RNIG894[15]\ : MX2C
      port map(A => \addr_data_vector[47]\, B => 
        addr_data_vector_79, S => sel_data_0(1), Y => N_1284);
    
    \update_r[1]\ : DFN1C0
      port map(D => update_and_sel_5(3), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \update_r[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_17\ : OR2A
      port map(A => nb_burst_available(7), B => 
        \un2_nb_send_next[7]\, Y => N_28);
    
    \FSM_SELECT_ADDRESS.state7_0_I_43\ : AO1A
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), C => nb_burst_available(5), Y => 
        \ACT_LT2_E[2]\);
    
    \update_r_RNI1KV4_0[0]\ : OR2
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => \un1_state_12_3_0[4]\);
    
    un1_address_m57 : AX1C
      port map(A => \addr_data_vector[52]\, B => N_34_0, C => 
        \addr_data_vector[53]\, Y => \un1_address[21]\);
    
    un1_address_m20_m7_i_1 : NOR2B
      port map(A => \addr_data_vector[40]\, B => 
        \addr_data_vector[41]\, Y => m20_m7_i_1);
    
    un2_nb_send_next_I_8 : NOR2B
      port map(A => \nb_send[1]_net_1\, B => \nb_send[0]_net_1\, 
        Y => N_38);
    
    un1_address_m40_m6_0_a2 : NOR3A
      port map(A => m40_m6_0_a2_6, B => m36_m6_0_a2_4_i, C => 
        N_13_0, Y => N_41);
    
    \FSM_SELECT_ADDRESS.state7_0_I_23\ : AO1C
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), C => N_28, Y => N_34);
    
    \FSM_SELECT_ADDRESS.state7_0_I_26\ : OA1A
      port map(A => N_32, B => N_34, C => N_33, Y => N_37);
    
    \address_RNO[22]\ : MX2
      port map(A => \un1_address[22]\, B => addr_data_f1(22), S
         => \state[0]_net_1\, Y => \address_7[22]\);
    
    un2_nb_send_next_I_27 : AND2
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        Y => \DWACT_FINC_E[1]\);
    
    un1_address_m49 : XOR2
      port map(A => N_2, B => \addr_data_vector[35]\, Y => 
        N_50_i_0);
    
    \address_RNIQNMA[3]\ : MX2C
      port map(A => \addr_data_vector[35]\, B => 
        addr_data_vector_67, S => sel_data_0(1), Y => N_1300);
    
    \address[9]\ : DFN1C0
      port map(D => \address_7[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[41]\);
    
    \address_RNO[18]\ : MX2
      port map(A => \un1_address[18]\, B => addr_data_f1(18), S
         => \state[0]_net_1\, Y => \address_7[18]\);
    
    \address_RNIKVLA[0]\ : MX2C
      port map(A => \addr_data_vector[32]\, B => 
        addr_data_vector_64, S => sel_data_0(1), Y => N_1297);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \address_RNI8894[11]\ : MX2C
      port map(A => \addr_data_vector[43]\, B => 
        addr_data_vector_75, S => sel_data_0(1), Y => N_1294);
    
    \address_RNO[7]\ : MX2
      port map(A => N_1_i_0, B => addr_data_f1(7), S => 
        \state_0[0]_net_1\, Y => \address_7[7]\);
    
    \address[6]\ : DFN1C0
      port map(D => \address_7[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[38]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_59\ : OR2A
      port map(A => \un2_nb_send_next[3]\, B => 
        nb_burst_available(3), Y => \ACT_LT4_E[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_1\ : XNOR2
      port map(A => \un2_nb_send_next[10]\, B => 
        nb_burst_available(10), Y => \DWACT_BL_EQUAL_0_E[4]\);
    
    un1_address_m23 : NOR3C
      port map(A => \addr_data_vector[44]\, B => m20_N_17_i_0, C
         => \addr_data_vector[45]\, Y => N_24_0);
    
    status_full_err_RNO : AO1
      port map(A => \state[2]_net_1\, B => N_129, C => 
        un1_state_5_i_0, Y => N_110);
    
    \state_0[0]\ : DFN1C0
      port map(D => N_118, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state_0[0]_net_1\);
    
    \address_RNO[8]\ : MX2
      port map(A => N_15_0_i_0, B => addr_data_f1(8), S => 
        \state_0[0]_net_1\, Y => \address_7[8]\);
    
    un2_nb_send_next_I_52 : XOR2
      port map(A => N_7, B => \nb_send[9]_net_1\, Y => 
        \un2_nb_send_next[9]\);
    
    \address_RNIC894[13]\ : MX2C
      port map(A => \addr_data_vector[45]\, B => 
        addr_data_vector_77, S => sel_data_0(1), Y => N_1282);
    
    \address[11]\ : DFN1C0
      port map(D => \address_7[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[43]\);
    
    un1_address_m20_m3_e : OR2B
      port map(A => m20_m3_e_0, B => N_69, Y => m20_m3_e);
    
    \address[31]\ : DFN1C0
      port map(D => \address_7[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[63]\);
    
    un1_address_m36_m6_0_a2_4_6 : NOR3C
      port map(A => \addr_data_vector[51]\, B => 
        \addr_data_vector[50]\, C => m36_m6_0_a2_4_4, Y => 
        m36_m6_0_a2_4_6);
    
    \FSM_SELECT_ADDRESS.state7_0_I_55\ : OR2A
      port map(A => nb_burst_available(2), B => 
        \un2_nb_send_next[2]\, Y => \ACT_LT4_E[4]\);
    
    un1_address_m56 : XOR2
      port map(A => N_31_0, B => \addr_data_vector[50]\, Y => 
        \un1_address[18]\);
    
    \address_RNO[2]\ : MX2
      port map(A => N_40_i_0, B => addr_data_f1(2), S => 
        \state_0[0]_net_1\, Y => \address_7[2]\);
    
    un1_address_m44 : OR3B
      port map(A => \addr_data_vector[58]\, B => 
        \addr_data_vector[59]\, C => N_43, Y => N_45);
    
    \address_RNIOFMA[2]\ : MX2C
      port map(A => \addr_data_vector[34]\, B => 
        addr_data_vector_66, S => sel_data_0(1), Y => N_1299);
    
    \address_RNO[4]\ : MX2
      port map(A => N_51_i_0, B => addr_data_f1(4), S => 
        \state_0[0]_net_1\, Y => \address_7[4]\);
    
    un2_nb_send_next_I_19 : NOR2B
      port map(A => \nb_send[3]_net_1\, B => \DWACT_FINC_E[0]\, Y
         => N_30);
    
    \address_RNO[25]\ : MX2
      port map(A => \un1_address[25]\, B => addr_data_f1(25), S
         => \state[0]_net_1\, Y => \address_7[25]\);
    
    \address[21]\ : DFN1C0
      port map(D => \address_7[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[53]\);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    un1_address_m62 : AX1
      port map(A => N_43, B => \addr_data_vector[58]\, C => 
        \addr_data_vector[59]\, Y => \un1_address[27]\);
    
    un1_address_m32 : AX1C
      port map(A => \addr_data_vector[50]\, B => N_31_0, C => 
        \addr_data_vector[51]\, Y => \un1_address[19]\);
    
    un1_address_m12_e : OR3C
      port map(A => \addr_data_vector[36]\, B => N_69, C => 
        \addr_data_vector[37]\, Y => N_5_0);
    
    \address_RNO_5[31]\ : NOR2B
      port map(A => \addr_data_vector[58]\, B => 
        \addr_data_vector[59]\, Y => address_7_31_m6_e_1);
    
    un2_nb_send_next_I_9 : XOR2
      port map(A => N_38, B => \nb_send[2]_net_1\, Y => 
        \un2_nb_send_next[2]\);
    
    \state[1]\ : DFN1C0
      port map(D => N_116, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \state[1]_net_1\);
    
    \address_RNIF245[23]\ : MX2C
      port map(A => \addr_data_vector[55]\, B => 
        addr_data_vector_87, S => sel_data(1), Y => N_906);
    
    \address[17]\ : DFN1C0
      port map(D => \address_7[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[49]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_52\ : OR2A
      port map(A => nb_burst_available(1), B => 
        \un2_nb_send_next[1]\, Y => \ACT_LT4_E[1]\);
    
    \state_RNI40SU8_0[3]\ : OR2B
      port map(A => address_0_sqmuxa_0, B => state7, Y => 
        address_0_sqmuxa);
    
    un1_address_m65 : AX1C
      port map(A => \addr_data_vector[61]\, B => N_46, C => 
        \addr_data_vector[62]\, Y => \un1_address[30]\);
    
    un1_address_m52 : XNOR2
      port map(A => N_13_0, B => \addr_data_vector[39]\, Y => 
        N_1_i_0);
    
    \address[27]\ : DFN1C0
      port map(D => \address_7[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[59]\);
    
    \state_RNO[3]\ : NOR2A
      port map(A => \state[4]_net_1\, B => N_129, Y => N_113);
    
    un1_address_m21 : XOR2
      port map(A => m20_N_17_i_0, B => \addr_data_vector[44]\, Y
         => N_22_0_i_0);
    
    un1_address_m20_m7_i_3 : NOR3C
      port map(A => m20_m7_i_0, B => \addr_data_vector[42]\, C
         => m20_m7_i_1, Y => m20_m7_i_3);
    
    \nb_send_RNO[4]\ : NOR2B
      port map(A => \un2_nb_send_next[4]\, B => state7, Y => 
        \nb_send_5[4]\);
    
    \nb_send_RNO[10]\ : NOR2B
      port map(A => \un2_nb_send_next[10]\, B => state7, Y => 
        \nb_send_5[10]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_18\ : OR2A
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => N_29);
    
    un1_address_m55 : XOR2
      port map(A => N_24_0, B => \addr_data_vector[46]\, Y => 
        N_56_0_i_0);
    
    \address_RNO[31]\ : MX2C
      port map(A => \address_RNO_0[31]_net_1\, B => 
        \address_RNO_1[31]_net_1\, S => \address_RNO_2[31]_net_1\, 
        Y => \address_7[31]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_61\ : AOI1A
      port map(A => \ACT_LT4_E[3]\, B => \ACT_LT4_E[6]\, C => 
        \ACT_LT4_E[10]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\);
    
    un1_address_m20_m7_i_o5 : OR2A
      port map(A => \addr_data_vector[38]\, B => address_0_sqmuxa, 
        Y => m20_m7_i_o5);
    
    un1_address_m10_e : NOR2B
      port map(A => N_2, B => \addr_data_vector[35]\, Y => N_69);
    
    \FSM_SELECT_ADDRESS.state7_0_I_34\ : XNOR2
      port map(A => \un2_nb_send_next[4]\, B => 
        nb_burst_available(4), Y => \DWACT_BL_EQUAL_0_E[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_6\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E_0[0]\, B => 
        \DWACT_BL_EQUAL_0_E_0[1]\, C => \DWACT_BL_EQUAL_0_E[2]\, 
        Y => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\);
    
    \address_RNO[12]\ : MX2
      port map(A => N_22_0_i_0, B => addr_data_f1(12), S => 
        \state_0[0]_net_1\, Y => \address_7[12]\);
    
    un2_nb_send_next_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \nb_send[6]_net_1\, Y => N_17);
    
    \address_RNIK894[17]\ : MX2C
      port map(A => \addr_data_vector[49]\, B => 
        addr_data_vector_81, S => sel_data_0(1), Y => N_1286);
    
    un2_nb_send_next_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_12);
    
    \state_RNIEABE[1]\ : NOR2A
      port map(A => status_full_ack(1), B => N_131, Y => N_118);
    
    \FSM_SELECT_ADDRESS.state7_0_I_3\ : XNOR2
      port map(A => \un2_nb_send_next[8]\, B => 
        nb_burst_available(8), Y => \DWACT_BL_EQUAL_0_E[2]\);
    
    status_full_RNO : AO1A
      port map(A => state7, B => \state[3]_net_1\, C => 
        \state[2]_net_1\, Y => un1_state_11);
    
    \address[1]\ : DFN1E1C0
      port map(D => addr_data_f1(1), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        \addr_data_vector[33]\);
    
    \status_full\ : DFN1E1C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_11, Q => status_full(1));
    
    \update_r_RNI1KV4[0]\ : OR2B
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => un3_update_r);
    
    un1_address_m63 : XNOR2
      port map(A => N_45, B => \addr_data_vector[60]\, Y => 
        \un1_address[28]\);
    
    un1_address_m33 : NOR3C
      port map(A => \addr_data_vector[50]\, B => N_31_0, C => 
        \addr_data_vector[51]\, Y => N_34_0);
    
    un2_nb_send_next_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    \address_RNID245[22]\ : MX2C
      port map(A => \addr_data_vector[54]\, B => 
        addr_data_vector_86, S => sel_data(1), Y => N_905);
    
    \address_RNIM7MA[1]\ : MX2C
      port map(A => \addr_data_vector[33]\, B => 
        addr_data_vector_65, S => sel_data_0(1), Y => N_1298);
    
    \address_RNO[20]\ : MX2
      port map(A => \un1_address[20]\, B => addr_data_f1(20), S
         => \state[0]_net_1\, Y => \address_7[20]\);
    
    \nb_send[8]\ : DFN1E0C0
      port map(D => \nb_send_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[8]_net_1\);
    
    un1_address_m53 : XOR2
      port map(A => N_18_0, B => \addr_data_vector[42]\, Y => 
        N_54_0_i_0);
    
    un1_address_m40_m6_0_a2_0 : NOR2B
      port map(A => \addr_data_vector[55]\, B => 
        \addr_data_vector[43]\, Y => m40_m6_0_a2_0);
    
    un1_address_m40_m6_0_a2_1 : NOR2B
      port map(A => \addr_data_vector[44]\, B => 
        \addr_data_vector[54]\, Y => m40_m6_0_a2_1);
    
    \address_RNO_3[31]\ : NOR3C
      port map(A => \addr_data_vector[57]\, B => 
        \addr_data_vector[62]\, C => address_7_31_m6_e_1, Y => 
        address_7_31_m6_e_3);
    
    \state_RNI14MB[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => un3_update_r, Y => 
        address_0_sqmuxa_0);
    
    \nb_send[1]\ : DFN1E0C0
      port map(D => \nb_send_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_60\ : AOI1A
      port map(A => \ACT_LT4_E[7]\, B => \ACT_LT4_E[8]\, C => 
        \ACT_LT4_E[5]\, Y => \ACT_LT4_E[10]\);
    
    \state_RNO_1[4]\ : OR3A
      port map(A => \state_0[0]_net_1\, B => \state[3]_net_1\, C
         => \state[2]_net_1\, Y => N_124);
    
    \address_RNO[15]\ : MX2
      port map(A => N_26_0_i_0, B => addr_data_f1(15), S => 
        \state_0[0]_net_1\, Y => \address_7[15]\);
    
    un1_address_m20_m7_i : AOI1B
      port map(A => m20_m7_i_o5, B => m20_m3_e, C => m20_m7_i_4, 
        Y => m20_N_17_i_0);
    
    un2_nb_send_next_I_20 : XOR2
      port map(A => N_30, B => \nb_send[4]_net_1\, Y => 
        \un2_nb_send_next[4]\);
    
    un1_address_m42 : OR3C
      port map(A => \addr_data_vector[56]\, B => N_41, C => 
        \addr_data_vector[57]\, Y => N_43);
    
    \FSM_SELECT_ADDRESS.state7_0_I_68\ : AO1
      port map(A => \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, B => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, C => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, Y => 
        \DWACT_COMP0_E[2]\);
    
    \address_RNIN245[27]\ : MX2C
      port map(A => \addr_data_vector[59]\, B => 
        addr_data_vector_91, S => sel_data(1), Y => N_910);
    
    un2_nb_send_next_I_16 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_dma_send_1word is

    port( Lock             : out   std_logic;
          Request          : out   std_logic;
          HRESETn_c        : in    std_logic;
          HCLK_c           : in    std_logic;
          un1_time_send_ok : out   std_logic;
          time_select      : in    std_logic;
          Store            : in    std_logic;
          N_1012           : out   std_logic;
          Ready            : in    std_logic;
          Fault            : in    std_logic;
          time_send        : in    std_logic;
          Grant            : in    std_logic
        );

end lpp_dma_send_1word;

architecture DEF_ARCH of lpp_dma_send_1word is 

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un1_state_4_i_0, \state[1]_net_1\, \state[3]_net_1\, 
        \state_ns_i_a4_0[0]\, \state[0]_net_1\, \state[2]_net_1\, 
        un1_state_2, N_69, \state[4]_net_1\, N_66, N_58, N_60, 
        \state_ns[1]\, Request_4, N_61, Store_0, \state_ns[2]\, 
        \state_RNO[4]_net_1\, time_send_ok, time_send_ko, 
        \state_ns[3]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \state_RNI4AM7[1]\ : OR2
      port map(A => \state[1]_net_1\, B => \state[3]_net_1\, Y
         => un1_state_4_i_0);
    
    \state[1]\ : DFN1C0
      port map(D => \state_ns[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[1]_net_1\);
    
    \state_RNIFCT8[4]\ : NOR2B
      port map(A => time_send, B => \state[4]_net_1\, Y => 
        Request_4);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \state_RNIAJH31[3]\ : NOR2B
      port map(A => \state[3]_net_1\, B => Grant, Y => N_66);
    
    \state_RNI6OUR[2]\ : NOR2A
      port map(A => \state[2]_net_1\, B => N_61, Y => N_69);
    
    un1_state_2_0_o3 : NOR2A
      port map(A => Fault, B => Ready, Y => N_61);
    
    \state[4]\ : DFN1P0
      port map(D => \state_RNO[4]_net_1\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[4]_net_1\);
    
    \DMAIn.Request\ : DFN1E1C0
      port map(D => Request_4, CLK => HCLK_c, CLR => HRESETn_c, E
         => un1_state_2, Q => Request);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \state_RNO[4]\ : OA1C
      port map(A => time_send, B => \state_ns_i_a4_0[0]\, C => 
        N_58, Y => \state_RNO[4]_net_1\);
    
    \state_RNIKGB32[4]\ : OR3
      port map(A => N_69, B => \state[4]_net_1\, C => N_66, Y => 
        un1_state_2);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    send_ok : DFN1E0C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_58, Q => time_send_ok);
    
    \state_RNO[1]\ : NOR2A
      port map(A => \state[2]_net_1\, B => Fault, Y => 
        \state_ns[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DMAIn.Store_RNIVI9A\ : MX2
      port map(A => Store, B => Store_0, S => time_select, Y => 
        N_1012);
    
    \state_RNO_0[4]\ : OR2
      port map(A => \state[0]_net_1\, B => \state[2]_net_1\, Y
         => \state_ns_i_a4_0[0]\);
    
    \DMAIn.Store\ : DFN1E1C0
      port map(D => \state[4]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_2, Q => Store_0);
    
    \DMAIn.Lock\ : DFN1E1C0
      port map(D => time_send, CLK => HCLK_c, CLR => HRESETn_c, E
         => \state[4]_net_1\, Q => Lock);
    
    \state_RNO[2]\ : AO1
      port map(A => \state[2]_net_1\, B => N_61, C => N_66, Y => 
        \state_ns[2]\);
    
    \state_ns_i_o3[0]\ : NOR2B
      port map(A => Ready, B => Fault, Y => N_60);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \state_RNO[3]\ : AO1A
      port map(A => Grant, B => \state[3]_net_1\, C => Request_4, 
        Y => \state_ns[1]\);
    
    send_ko_RNI8BV9 : OR2
      port map(A => time_send_ok, B => time_send_ko, Y => 
        un1_time_send_ok);
    
    send_ko : DFN1E0C0
      port map(D => \state[0]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_58, Q => time_send_ko);
    
    \state[0]\ : DFN1C0
      port map(D => \state[1]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[0]_net_1\);
    
    \state_RNIA2L31[2]\ : AO1A
      port map(A => N_60, B => \state[2]_net_1\, C => 
        un1_state_4_i_0, Y => N_58);
    
    \state[3]\ : DFN1C0
      port map(D => \state_ns[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\ is

    port( nb_burst_available  : in    std_logic_vector(10 downto 0);
          status_full_err     : out   std_logic_vector(3 to 3);
          status_full         : out   std_logic_vector(3 to 3);
          sel_data            : in    std_logic_vector(1 to 1);
          sel_data_0          : in    std_logic_vector(1 to 1);
          update_and_sel_1    : in    std_logic_vector(7 downto 6);
          addr_data_f3        : in    std_logic_vector(31 downto 0);
          status_full_ack     : in    std_logic_vector(3 to 3);
          addr_data_vector_61 : out   std_logic;
          addr_data_vector_60 : out   std_logic;
          addr_data_vector_27 : in    std_logic;
          addr_data_vector_25 : in    std_logic;
          addr_data_vector_24 : in    std_logic;
          addr_data_vector_22 : in    std_logic;
          addr_data_vector_20 : in    std_logic;
          addr_data_vector_0  : in    std_logic;
          addr_data_vector_6  : in    std_logic;
          addr_data_vector_4  : in    std_logic;
          addr_data_vector_3  : in    std_logic;
          addr_data_vector_2  : in    std_logic;
          addr_data_vector_1  : in    std_logic;
          addr_data_vector_14 : in    std_logic;
          addr_data_vector_12 : in    std_logic;
          addr_data_vector_10 : in    std_logic;
          addr_data_vector_8  : in    std_logic;
          addr_data_vector_63 : out   std_logic;
          addr_data_vector_90 : out   std_logic;
          addr_data_vector_87 : out   std_logic;
          addr_data_vector_85 : out   std_logic;
          addr_data_vector_62 : out   std_logic;
          addr_data_vector_69 : out   std_logic;
          addr_data_vector_73 : out   std_logic;
          addr_data_vector_71 : out   std_logic;
          addr_data_vector_77 : out   std_logic;
          addr_data_vector_79 : out   std_logic;
          addr_data_vector_82 : out   std_logic;
          addr_data_vector_83 : out   std_logic;
          addr_data_vector_75 : out   std_logic;
          addr_data_vector_80 : out   std_logic;
          addr_data_vector_81 : out   std_logic;
          N_914               : out   std_logic;
          N_912               : out   std_logic;
          N_911               : out   std_logic;
          N_909               : out   std_logic;
          N_907               : out   std_logic;
          N_1301              : out   std_logic;
          N_1293              : out   std_logic;
          N_1291              : out   std_logic;
          N_1290              : out   std_logic;
          N_1289              : out   std_logic;
          N_1288              : out   std_logic;
          N_1287              : out   std_logic;
          N_1285              : out   std_logic;
          N_1283              : out   std_logic;
          N_1281              : out   std_logic;
          HRESETn_c           : in    std_logic;
          HCLK_c              : in    std_logic
        );

end 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\;

architecture DEF_ARCH of 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\ is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \state_0[0]_net_1\, \state_RNIKABE[1]_net_1\, N_38, 
        \nb_send[1]_net_1\, \nb_send[0]_net_1\, N_30, 
        \nb_send[3]_net_1\, \DWACT_FINC_E[0]\, N_7, 
        \nb_send[8]_net_1\, \DWACT_FINC_E[4]\, m40_m6_0_a2_7, 
        m40_m6_0_a2_2, m40_m6_0_a2_1, m40_m6_0_a2_6, 
        m40_m6_0_a2_4, \addr_data_vector[114]\, 
        \addr_data_vector[112]\, m24_m5_0_a2_5, 
        \addr_data_vector[106]\, m24_m5_0_a2_3, m24_m5_0_a2_4, 
        \addr_data_vector[103]\, \addr_data_vector[110]\, 
        m24_m5_0_a2_1, \addr_data_vector[108]\, 
        \addr_data_vector[104]\, \un1_state_12_3_0[4]\, 
        \update_r_i[0]\, \update_r[1]_net_1\, un1_state_5_i_0, 
        \state[4]_net_1\, \state[3]_net_1\, \state_ns_i_0[3]\, 
        N_131, \un1_state_12[4]\, \un1_state_12_2[4]\, 
        \un1_address[6]\, address_0_sqmuxa, 
        \addr_data_vector[102]\, N_5_0, \state_RNO[1]_net_1\, 
        N_129, \state[1]_net_1\, \state_ns[0]\, N_125, N_124, 
        N_110, \state[2]_net_1\, state7, un3_update_r, N_25_0_i_0, 
        N_13_0, N_15_0_i_0, N_16_0, N_17_0_i_0, 
        \addr_data_vector[105]\, N_19_0, N_20_0_i_0, 
        \addr_data_vector[107]\, N_22_0_i_0, N_23_0, N_26_0_i_0, 
        \addr_data_vector[111]\, N_28_0_i_0, N_29_0, N_30_0_i_0, 
        \addr_data_vector[113]\, N_32_0, N_33_0, 
        \addr_data_vector[115]\, N_35_0, \addr_data_vector[116]\, 
        N_36_0, N_37_0, \addr_data_vector[117]\, N_39, 
        \addr_data_vector[118]\, \addr_data_vector[119]\, 
        N_40_i_0, N_42, \addr_data_vector[120]\, N_44, 
        \addr_data_vector[122]\, N_46, \addr_data_vector[124]\, 
        N_47, \addr_data_vector[125]\, N_49_i_0, 
        \addr_data_vector[127]\, N_50_i_0, \addr_data_vector[98]\, 
        N_51_i_0, N_69, \addr_data_vector[100]\, N_52_i_0, 
        \addr_data_vector[101]\, N_1_i_0, N_54_0_i_0, N_55_0_i_0, 
        \addr_data_vector[109]\, N_57_0, N_58_0, N_59_0, N_60_0, 
        N_61_0, \addr_data_vector[121]\, N_62, N_63_0, 
        \addr_data_vector[123]\, N_64_0, N_65_0, N_66_0, 
        \addr_data_vector[126]\, \addr_data_vector[99]\, 
        \address_7[2]\, \address_7[3]\, \address_7[4]\, 
        \address_7[5]\, \address_7[6]\, \address_7[7]\, 
        \address_7[8]\, \address_7[9]\, \address_7[10]\, 
        \address_7[11]\, \address_7[12]\, \address_7[13]\, 
        \address_7[15]\, \address_7[16]\, \address_7[17]\, 
        \address_7[18]\, \address_7[19]\, \state[0]_net_1\, 
        \address_7[20]\, \address_7[21]\, \address_7[22]\, 
        \address_7[23]\, \address_7[24]\, \address_7[25]\, 
        \address_7[26]\, \address_7[27]\, \address_7[28]\, 
        \address_7[29]\, \address_7[30]\, \address_7[31]\, 
        N_56_0_i_0, un1_state_9, \nb_send_5[0]\, \nb_send_5[1]\, 
        I_5_19, \nb_send_5[2]\, I_9_19, \nb_send_5[3]\, I_13_19, 
        \nb_send_5[4]\, I_20_11, \nb_send_5[5]\, I_24_3, 
        \nb_send_5[6]\, I_31_4, \nb_send_5[7]\, I_38_3, 
        \nb_send_5[8]\, I_45_3, \nb_send_5[9]\, I_52_3, 
        \nb_send_5[10]\, I_56_3, N_127, \state_RNO_0[3]\, 
        \state_ns[2]\, un1_state_11, \address_7[14]\, 
        \nb_send[2]_net_1\, \nb_send[4]_net_1\, 
        \nb_send[5]_net_1\, \nb_send[6]_net_1\, 
        \nb_send[7]_net_1\, \nb_send[9]_net_1\, 
        \nb_send[10]_net_1\, N_4, \DWACT_FINC_E[2]\, 
        \DWACT_FINC_E[3]\, N_12, N_17, N_22, \DWACT_FINC_E[1]\, 
        N_27, N_35, \DWACT_COMP0_E[1]\, \DWACT_COMP0_E[2]\, 
        \DWACT_COMP0_E[0]\, \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, \ACT_LT4_E[3]\, 
        \ACT_LT4_E[6]\, \ACT_LT4_E[10]\, \ACT_LT4_E[7]\, 
        \ACT_LT4_E[8]\, \ACT_LT4_E[5]\, \ACT_LT4_E[4]\, 
        \ACT_LT4_E[0]\, \ACT_LT4_E[1]\, \ACT_LT4_E[2]\, 
        \ACT_LT2_E[0]\, \ACT_LT2_E[1]\, \ACT_LT2_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, N_37, 
        N_36, N_35_1, N_32, N_34, N_33, N_31, N_28, N_29, N_30_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, 
        \DWACT_BL_EQUAL_0_E[4]\, \DWACT_BL_EQUAL_0_E[3]\, 
        \DWACT_BL_EQUAL_0_E_0[0]\, \DWACT_BL_EQUAL_0_E_0[1]\, 
        \DWACT_BL_EQUAL_0_E[2]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    addr_data_vector_63 <= \addr_data_vector[99]\;
    addr_data_vector_90 <= \addr_data_vector[126]\;
    addr_data_vector_87 <= \addr_data_vector[123]\;
    addr_data_vector_85 <= \addr_data_vector[121]\;
    addr_data_vector_62 <= \addr_data_vector[98]\;
    addr_data_vector_69 <= \addr_data_vector[105]\;
    addr_data_vector_73 <= \addr_data_vector[109]\;
    addr_data_vector_71 <= \addr_data_vector[107]\;
    addr_data_vector_77 <= \addr_data_vector[113]\;
    addr_data_vector_79 <= \addr_data_vector[115]\;
    addr_data_vector_82 <= \addr_data_vector[118]\;
    addr_data_vector_83 <= \addr_data_vector[119]\;
    addr_data_vector_75 <= \addr_data_vector[111]\;
    addr_data_vector_80 <= \addr_data_vector[116]\;
    addr_data_vector_81 <= \addr_data_vector[117]\;

    \address[16]\ : DFN1C0
      port map(D => \address_7[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[112]\);
    
    \address[10]\ : DFN1C0
      port map(D => \address_7[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[106]\);
    
    \state[0]\ : DFN1C0
      port map(D => \state_RNIKABE[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state[0]_net_1\);
    
    \address[30]\ : DFN1C0
      port map(D => \address_7[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[126]\);
    
    un1_address_m45 : OR3B
      port map(A => \addr_data_vector[123]\, B => 
        \addr_data_vector[124]\, C => N_44, Y => N_46);
    
    \address_RNO[26]\ : MX2
      port map(A => N_62, B => addr_data_f3(26), S => 
        \state[0]_net_1\, Y => \address_7[26]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_25\ : AO1C
      port map(A => I_52_3, B => nb_burst_available(9), C => N_31, 
        Y => N_36);
    
    un1_address_m61 : AX1
      port map(A => N_42, B => \addr_data_vector[121]\, C => 
        \addr_data_vector[122]\, Y => N_62);
    
    un1_address_m31 : OR3B
      port map(A => \addr_data_vector[113]\, B => 
        \addr_data_vector[114]\, C => N_29_0, Y => N_32_0);
    
    \address[26]\ : DFN1C0
      port map(D => \address_7[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[122]\);
    
    \address[20]\ : DFN1C0
      port map(D => \address_7[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[116]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_42\ : AO1C
      port map(A => I_20_11, B => nb_burst_available(4), C => 
        I_24_3, Y => \ACT_LT2_E[1]\);
    
    \state_RNO_0[2]\ : NOR3B
      port map(A => N_129, B => \state[2]_net_1\, C => 
        status_full_ack(3), Y => N_127);
    
    \FSM_SELECT_ADDRESS.state7_0_I_57\ : NOR2A
      port map(A => \ACT_LT4_E[4]\, B => \ACT_LT4_E[5]\, Y => 
        \ACT_LT4_E[6]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_36\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[1]\, B => 
        \DWACT_BL_EQUAL_0_E[0]\, Y => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\);
    
    un1_address_m51 : AX1C
      port map(A => \addr_data_vector[100]\, B => N_69, C => 
        \addr_data_vector[101]\, Y => N_52_i_0);
    
    \address[12]\ : DFN1C0
      port map(D => \address_7[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[108]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_22\ : OA1A
      port map(A => I_52_3, B => nb_burst_available(9), C => N_29, 
        Y => N_33);
    
    \address_RNO[29]\ : MX2
      port map(A => N_65_0, B => addr_data_f3(29), S => 
        \state[0]_net_1\, Y => \address_7[29]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_8\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\, B => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\, Y => 
        \DWACT_COMP0_E[1]\);
    
    un1_address_m19 : XOR2
      port map(A => N_19_0, B => \addr_data_vector[107]\, Y => 
        N_20_0_i_0);
    
    \address[22]\ : DFN1C0
      port map(D => \address_7[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[118]\);
    
    \address_RNO[23]\ : MX2
      port map(A => N_39, B => addr_data_f3(23), S => 
        \state[0]_net_1\, Y => \address_7[23]\);
    
    \address[2]\ : DFN1C0
      port map(D => \address_7[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[98]\);
    
    un2_nb_send_next_I_13 : XOR2
      port map(A => N_35, B => \nb_send[3]_net_1\, Y => I_13_19);
    
    un1_address_m43 : OR3B
      port map(A => \addr_data_vector[121]\, B => 
        \addr_data_vector[122]\, C => N_42, Y => N_44);
    
    \FSM_SELECT_ADDRESS.state7_0_I_54\ : AOI1A
      port map(A => \ACT_LT4_E[0]\, B => \ACT_LT4_E[1]\, C => 
        \ACT_LT4_E[2]\, Y => \ACT_LT4_E[3]\);
    
    \address_RNO[24]\ : MX2
      port map(A => N_60_0, B => addr_data_f3(24), S => 
        \state[0]_net_1\, Y => \address_7[24]\);
    
    \address_RNO[10]\ : MX2
      port map(A => N_54_0_i_0, B => addr_data_f3(10), S => 
        \state_0[0]_net_1\, Y => \address_7[10]\);
    
    \status_full_err\ : DFN1E0C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_110, Q => status_full_err(3));
    
    un2_nb_send_next_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \nb_send[8]_net_1\, C
         => \nb_send[9]_net_1\, Y => N_4);
    
    un1_address_m18 : NOR3C
      port map(A => \addr_data_vector[105]\, B => N_16_0, C => 
        \addr_data_vector[106]\, Y => N_19_0);
    
    \nb_send_RNO[1]\ : NOR2B
      port map(A => I_5_19, B => state7, Y => \nb_send_5[1]\);
    
    \address_RNIA894[12]\ : MX2C
      port map(A => addr_data_vector_8, B => 
        \addr_data_vector[108]\, S => sel_data_0(1), Y => N_1281);
    
    \address_RNI40OA[8]\ : MX2C
      port map(A => addr_data_vector_4, B => 
        \addr_data_vector[104]\, S => sel_data_0(1), Y => N_1291);
    
    \FSM_SELECT_ADDRESS.state7_0_I_51\ : NOR2B
      port map(A => \nb_send[0]_net_1\, B => 
        nb_burst_available(0), Y => \ACT_LT4_E[0]\);
    
    un2_nb_send_next_I_31 : XOR2
      port map(A => N_22, B => \nb_send[6]_net_1\, Y => I_31_4);
    
    \nb_send[9]\ : DFN1E0C0
      port map(D => \nb_send_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[9]_net_1\);
    
    \address_RNO[9]\ : MX2
      port map(A => N_17_0_i_0, B => addr_data_f3(9), S => 
        \state_0[0]_net_1\, Y => \address_7[9]\);
    
    \address[5]\ : DFN1C0
      port map(D => \address_7[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[101]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_5\ : XNOR2
      port map(A => I_38_3, B => nb_burst_available(7), Y => 
        \DWACT_BL_EQUAL_0_E_0[1]\);
    
    \address[15]\ : DFN1C0
      port map(D => \address_7[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[111]\);
    
    \address[13]\ : DFN1C0
      port map(D => \address_7[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[109]\);
    
    \update_r_RNI5KV4[0]\ : OR2B
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => un3_update_r);
    
    \state[4]\ : DFN1P0
      port map(D => \state_ns[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[4]_net_1\);
    
    \nb_send_RNO[9]\ : NOR2B
      port map(A => I_52_3, B => state7, Y => \nb_send_5[9]\);
    
    \address[19]\ : DFN1C0
      port map(D => \address_7[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[115]\);
    
    \address_RNII894[16]\ : MX2C
      port map(A => addr_data_vector_12, B => 
        \addr_data_vector[112]\, S => sel_data_0(1), Y => N_1285);
    
    \address[25]\ : DFN1C0
      port map(D => \address_7[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[121]\);
    
    un2_nb_send_next_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => \nb_send[5]_net_1\, Y => N_22);
    
    \address_RNIL245[26]\ : MX2C
      port map(A => addr_data_vector_22, B => 
        \addr_data_vector[122]\, S => sel_data(1), Y => N_909);
    
    \address[23]\ : DFN1C0
      port map(D => \address_7[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[119]\);
    
    un1_address_m14 : AX1C
      port map(A => \addr_data_vector[103]\, B => N_13_0, C => 
        \addr_data_vector[104]\, Y => N_15_0_i_0);
    
    un1_address_m29 : XNOR2
      port map(A => N_29_0, B => \addr_data_vector[113]\, Y => 
        N_30_0_i_0);
    
    un2_nb_send_next_I_12 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => N_35);
    
    \FSM_SELECT_ADDRESS.state7_0_I_19\ : NOR2A
      port map(A => nb_burst_available(6), B => I_31_4, Y => 
        N_30_0);
    
    \address_RNIH245[24]\ : MX2C
      port map(A => addr_data_vector_20, B => 
        \addr_data_vector[120]\, S => sel_data(1), Y => N_907);
    
    \state_RNIKABE[1]\ : NOR2A
      port map(A => status_full_ack(3), B => N_131, Y => 
        \state_RNIKABE[1]_net_1\);
    
    \address[29]\ : DFN1C0
      port map(D => \address_7[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[125]\);
    
    \address[18]\ : DFN1C0
      port map(D => \address_7[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[114]\);
    
    \nb_send_RNO[6]\ : NOR2B
      port map(A => I_31_4, B => state7, Y => \nb_send_5[6]\);
    
    \address_RNO[21]\ : MX2
      port map(A => N_58_0, B => addr_data_f3(21), S => 
        \state[0]_net_1\, Y => \address_7[21]\);
    
    \address_RNO[16]\ : MX2
      port map(A => N_28_0_i_0, B => addr_data_f3(16), S => 
        \state_0[0]_net_1\, Y => \address_7[16]\);
    
    un2_nb_send_next_I_51 : NOR2B
      port map(A => \nb_send[8]_net_1\, B => \DWACT_FINC_E[4]\, Y
         => N_7);
    
    \address[0]\ : DFN1E1C0
      port map(D => addr_data_f3(0), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        addr_data_vector_60);
    
    un1_address_m28 : OR3B
      port map(A => \addr_data_vector[111]\, B => 
        \addr_data_vector[112]\, C => N_25_0_i_0, Y => N_29_0);
    
    status_full_err_RNO_0 : OR2
      port map(A => \state[4]_net_1\, B => \state[3]_net_1\, Y
         => un1_state_5_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_address_m41 : OR3B
      port map(A => m40_m6_0_a2_7, B => \addr_data_vector[120]\, 
        C => N_25_0_i_0, Y => N_42);
    
    \address_RNO[27]\ : MX2
      port map(A => N_63_0, B => addr_data_f3(27), S => 
        \state[0]_net_1\, Y => \address_7[27]\);
    
    \address[4]\ : DFN1C0
      port map(D => \address_7[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[100]\);
    
    \address[28]\ : DFN1C0
      port map(D => \address_7[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[124]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_7\ : AND2
      port map(A => \DWACT_BL_EQUAL_0_E[4]\, B => 
        \DWACT_BL_EQUAL_0_E[3]\, Y => 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1]\);
    
    \nb_send_RNO[2]\ : NOR2B
      port map(A => I_9_19, B => state7, Y => \nb_send_5[2]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \state_RNO_0[4]\ : OR3B
      port map(A => N_131, B => N_129, C => \state[3]_net_1\, Y
         => N_125);
    
    \address_RNI6894[10]\ : MX2C
      port map(A => addr_data_vector_6, B => 
        \addr_data_vector[106]\, S => sel_data_0(1), Y => N_1293);
    
    \FSM_SELECT_ADDRESS.state7_0_I_58\ : NOR2A
      port map(A => I_9_19, B => nb_burst_available(2), Y => 
        \ACT_LT4_E[7]\);
    
    \nb_send_RNO[7]\ : NOR2B
      port map(A => I_38_3, B => state7, Y => \nb_send_5[7]\);
    
    un2_nb_send_next_I_24 : XOR2
      port map(A => N_27, B => \nb_send[5]_net_1\, Y => I_24_3);
    
    un2_nb_send_next_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \nb_send[3]_net_1\, C
         => \nb_send[4]_net_1\, Y => N_27);
    
    un1_address_ADD_32x32_fast_I164_Y_0 : XNOR3
      port map(A => address_0_sqmuxa, B => 
        \addr_data_vector[102]\, C => N_5_0, Y => 
        \un1_address[6]\);
    
    \address_RNO[19]\ : MX2
      port map(A => N_33_0, B => addr_data_f3(19), S => 
        \state[0]_net_1\, Y => \address_7[19]\);
    
    \nb_send[7]\ : DFN1E0C0
      port map(D => \nb_send_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[7]_net_1\);
    
    \address_RNO[13]\ : MX2
      port map(A => N_55_0_i_0, B => addr_data_f3(13), S => 
        \state_0[0]_net_1\, Y => \address_7[13]\);
    
    \address[14]\ : DFN1C0
      port map(D => \address_7[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[110]\);
    
    \state_RNO[1]\ : OA1C
      port map(A => N_129, B => \state[1]_net_1\, C => 
        \state_ns_i_0[3]\, Y => \state_RNO[1]_net_1\);
    
    \nb_send[0]\ : DFN1E0C0
      port map(D => \nb_send_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[0]_net_1\);
    
    \state_RNILNSP8[3]\ : OR2B
      port map(A => \state[3]_net_1\, B => state7, Y => 
        \un1_state_12_2[4]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_53\ : AND2A
      port map(A => nb_burst_available(1), B => I_5_19, Y => 
        \ACT_LT4_E[2]\);
    
    un1_address_m40_m6_0_a2_4 : NOR3C
      port map(A => \addr_data_vector[111]\, B => 
        \addr_data_vector[119]\, C => \addr_data_vector[118]\, Y
         => m40_m6_0_a2_4);
    
    \nb_send[6]\ : DFN1E0C0
      port map(D => \nb_send_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[6]_net_1\);
    
    \nb_send[10]\ : DFN1E0C0
      port map(D => \nb_send_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[10]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_56\ : NOR2A
      port map(A => nb_burst_available(3), B => I_13_19, Y => 
        \ACT_LT4_E[5]\);
    
    \address_RNO[14]\ : MX2
      port map(A => N_56_0_i_0, B => addr_data_f3(14), S => 
        \state[0]_net_1\, Y => \address_7[14]\);
    
    \nb_send_RNO[3]\ : NOR2B
      port map(A => I_13_19, B => state7, Y => \nb_send_5[3]\);
    
    \nb_send[2]\ : DFN1E0C0
      port map(D => \nb_send_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[2]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_27\ : OA1
      port map(A => N_37, B => N_36, C => N_35_1, Y => 
        \DWACT_COMP0_E[0]\);
    
    \address[24]\ : DFN1C0
      port map(D => \address_7[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[120]\);
    
    un1_address_m27 : AX1
      port map(A => N_25_0_i_0, B => \addr_data_vector[111]\, C
         => \addr_data_vector[112]\, Y => N_28_0_i_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un1_address_m60 : XNOR2
      port map(A => N_42, B => \addr_data_vector[121]\, Y => 
        N_61_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_44\ : AND3A
      port map(A => \ACT_LT2_E[0]\, B => \ACT_LT2_E[1]\, C => 
        \ACT_LT2_E[2]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\);
    
    \nb_send[4]\ : DFN1E0C0
      port map(D => \nb_send_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[4]_net_1\);
    
    un1_address_m16 : XOR2
      port map(A => N_16_0, B => \addr_data_vector[105]\, Y => 
        N_17_0_i_0);
    
    un2_nb_send_next_I_45 : XOR2
      port map(A => N_12, B => \nb_send[8]_net_1\, Y => I_45_3);
    
    \nb_send_RNO[0]\ : NOR2A
      port map(A => state7, B => \nb_send[0]_net_1\, Y => 
        \nb_send_5[0]\);
    
    \nb_send_RNO[8]\ : NOR2B
      port map(A => I_45_3, B => state7, Y => \nb_send_5[8]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_41\ : AND2A
      port map(A => nb_burst_available(5), B => I_24_3, Y => 
        \ACT_LT2_E[0]\);
    
    \state_RNO[4]\ : OR3C
      port map(A => N_125, B => N_124, C => \un1_state_12_2[4]\, 
        Y => \state_ns[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_4\ : XNOR2
      port map(A => I_52_3, B => nb_burst_available(9), Y => 
        \DWACT_BL_EQUAL_0_E[3]\);
    
    \address[8]\ : DFN1C0
      port map(D => \address_7[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[104]\);
    
    un1_address_m40_m6_0_a2_2 : NOR2B
      port map(A => \addr_data_vector[114]\, B => 
        \addr_data_vector[115]\, Y => m40_m6_0_a2_2);
    
    un1_address_m50 : XOR2
      port map(A => N_69, B => \addr_data_vector[100]\, Y => 
        N_51_i_0);
    
    un1_address_m39 : XOR2
      port map(A => \un1_state_12[4]\, B => 
        \addr_data_vector[98]\, Y => N_40_i_0);
    
    \FSM_SELECT_ADDRESS.state7_0_I_24\ : OR2A
      port map(A => I_56_3, B => nb_burst_available(10), Y => 
        N_35_1);
    
    \state_ns_i_a2[1]\ : NOR2A
      port map(A => update_and_sel_1(6), B => update_and_sel_1(7), 
        Y => N_129);
    
    \address_RNO[6]\ : MX2
      port map(A => \un1_address[6]\, B => addr_data_f3(6), S => 
        \state_0[0]_net_1\, Y => \address_7[6]\);
    
    \update_r_RNIQBSU8[0]\ : NOR2
      port map(A => \un1_state_12_3_0[4]\, B => 
        \un1_state_12_2[4]\, Y => \un1_state_12[4]\);
    
    \state_RNO[2]\ : AO1A
      port map(A => state7, B => \state[3]_net_1\, C => N_127, Y
         => \state_ns[2]\);
    
    \address_RNO[28]\ : MX2
      port map(A => N_64_0, B => addr_data_f3(28), S => 
        \state[0]_net_1\, Y => \address_7[28]\);
    
    \address_RNO[11]\ : MX2
      port map(A => N_20_0_i_0, B => addr_data_f3(11), S => 
        \state_0[0]_net_1\, Y => \address_7[11]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_21\ : AO1C
      port map(A => nb_burst_available(7), B => I_38_3, C => 
        N_30_0, Y => N_32);
    
    \FSM_SELECT_ADDRESS.state7_0_I_73\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => state7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_35\ : XNOR2
      port map(A => I_24_3, B => nb_burst_available(5), Y => 
        \DWACT_BL_EQUAL_0_E[1]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_2\ : XNOR2
      port map(A => I_31_4, B => nb_burst_available(6), Y => 
        \DWACT_BL_EQUAL_0_E_0[0]\);
    
    un1_address_m38 : AX1C
      port map(A => \addr_data_vector[118]\, B => N_37_0, C => 
        \addr_data_vector[119]\, Y => N_39);
    
    un1_address_m12 : AO13
      port map(A => address_0_sqmuxa, B => 
        \addr_data_vector[102]\, C => N_5_0, Y => N_13_0);
    
    un1_address_m59 : AX1
      port map(A => N_25_0_i_0, B => m40_m6_0_a2_7, C => 
        \addr_data_vector[120]\, Y => N_60_0);
    
    \update_r[0]\ : DFN1P0
      port map(D => update_and_sel_1(6), CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \update_r_i[0]\);
    
    un2_nb_send_next_I_5 : XOR2
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        Y => I_5_19);
    
    un1_address_m40_m6_0_a2_6 : NOR3C
      port map(A => \addr_data_vector[117]\, B => 
        \addr_data_vector[116]\, C => m40_m6_0_a2_4, Y => 
        m40_m6_0_a2_6);
    
    \address_RNO[17]\ : MX2
      port map(A => N_30_0_i_0, B => addr_data_f3(17), S => 
        \state_0[0]_net_1\, Y => \address_7[17]\);
    
    \address_RNO[5]\ : MX2
      port map(A => N_52_i_0, B => addr_data_f3(5), S => 
        \state_0[0]_net_1\, Y => \address_7[5]\);
    
    un1_address_m15 : NOR3C
      port map(A => \addr_data_vector[103]\, B => N_13_0, C => 
        \addr_data_vector[104]\, Y => N_16_0);
    
    un1_address_m58 : XOR2
      port map(A => N_37_0, B => \addr_data_vector[118]\, Y => 
        N_59_0);
    
    \address_RNIU7NA[5]\ : MX2C
      port map(A => addr_data_vector_1, B => 
        \addr_data_vector[101]\, S => sel_data_0(1), Y => N_1288);
    
    un2_nb_send_next_I_56 : XOR2
      port map(A => N_4, B => \nb_send[10]_net_1\, Y => I_56_3);
    
    un2_nb_send_next_I_41 : AND2
      port map(A => \nb_send[6]_net_1\, B => \nb_send[7]_net_1\, 
        Y => \DWACT_FINC_E[3]\);
    
    \address_RNO[3]\ : MX2
      port map(A => N_50_i_0, B => addr_data_f3(3), S => 
        \state_0[0]_net_1\, Y => \address_7[3]\);
    
    \address[3]\ : DFN1C0
      port map(D => \address_7[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[99]\);
    
    \address_RNIR245[29]\ : MX2C
      port map(A => addr_data_vector_25, B => 
        \addr_data_vector[125]\, S => sel_data(1), Y => N_912);
    
    un2_nb_send_next_I_34 : AND3
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        C => \nb_send[5]_net_1\, Y => \DWACT_FINC_E[2]\);
    
    un1_address_m64 : XNOR2
      port map(A => N_46, B => \addr_data_vector[125]\, Y => 
        N_65_0);
    
    un1_address_m34 : AX1
      port map(A => N_32_0, B => \addr_data_vector[115]\, C => 
        \addr_data_vector[116]\, Y => N_35_0);
    
    \address_RNO[30]\ : MX2
      port map(A => N_66_0, B => addr_data_f3(30), S => 
        \state[0]_net_1\, Y => \address_7[30]\);
    
    \state_RNO_0[1]\ : OR2
      port map(A => status_full_ack(3), B => N_131, Y => 
        \state_ns_i_0[3]\);
    
    \nb_send[3]\ : DFN1E0C0
      port map(D => \nb_send_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[3]_net_1\);
    
    \state_RNIQBSU8_0[3]\ : AO1B
      port map(A => un3_update_r, B => state7, C => 
        \state[3]_net_1\, Y => un1_state_9);
    
    \FSM_SELECT_ADDRESS.state7_0_I_20\ : OR2A
      port map(A => nb_burst_available(10), B => I_56_3, Y => 
        N_31);
    
    un1_address_m54 : XOR2
      port map(A => N_23_0, B => \addr_data_vector[109]\, Y => 
        N_55_0_i_0);
    
    un1_address_m22 : NOR3C
      port map(A => \addr_data_vector[107]\, B => N_19_0, C => 
        \addr_data_vector[108]\, Y => N_23_0);
    
    \address[7]\ : DFN1C0
      port map(D => \address_7[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[103]\);
    
    un2_nb_send_next_I_38 : XOR2
      port map(A => N_17, B => \nb_send[7]_net_1\, Y => I_38_3);
    
    un1_address_m24_m5_0_a2_1 : NOR2B
      port map(A => \addr_data_vector[104]\, B => 
        \addr_data_vector[105]\, Y => m24_m5_0_a2_1);
    
    \nb_send[5]\ : DFN1E0C0
      port map(D => \nb_send_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[5]_net_1\);
    
    \nb_send_RNO[5]\ : NOR2B
      port map(A => I_24_3, B => state7, Y => \nb_send_5[5]\);
    
    un1_address_m25 : XNOR2
      port map(A => N_25_0_i_0, B => \addr_data_vector[111]\, Y
         => N_26_0_i_0);
    
    \state[3]\ : DFN1C0
      port map(D => \state_RNO_0[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    
    \update_r[1]\ : DFN1C0
      port map(D => update_and_sel_1(7), CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \update_r[1]_net_1\);
    
    un1_address_m40_m6_0_a2_7 : NOR3C
      port map(A => m40_m6_0_a2_2, B => m40_m6_0_a2_1, C => 
        m40_m6_0_a2_6, Y => m40_m6_0_a2_7);
    
    \FSM_SELECT_ADDRESS.state7_0_I_17\ : OR2A
      port map(A => nb_burst_available(7), B => I_38_3, Y => N_28);
    
    \FSM_SELECT_ADDRESS.state7_0_I_43\ : AO1A
      port map(A => I_20_11, B => nb_burst_available(4), C => 
        nb_burst_available(5), Y => \ACT_LT2_E[2]\);
    
    un1_address_m57 : XNOR2
      port map(A => N_36_0, B => \addr_data_vector[117]\, Y => 
        N_58_0);
    
    un2_nb_send_next_I_8 : NOR2B
      port map(A => \nb_send[1]_net_1\, B => \nb_send[0]_net_1\, 
        Y => N_38);
    
    \FSM_SELECT_ADDRESS.state7_0_I_23\ : AO1C
      port map(A => I_45_3, B => nb_burst_available(8), C => N_28, 
        Y => N_34);
    
    \FSM_SELECT_ADDRESS.state7_0_I_26\ : OA1A
      port map(A => N_32, B => N_34, C => N_33, Y => N_37);
    
    \address_RNI0GNA[6]\ : MX2C
      port map(A => addr_data_vector_2, B => 
        \addr_data_vector[102]\, S => sel_data_0(1), Y => N_1289);
    
    \address_RNO[22]\ : MX2
      port map(A => N_59_0, B => addr_data_f3(22), S => 
        \state[0]_net_1\, Y => \address_7[22]\);
    
    un2_nb_send_next_I_27 : AND2
      port map(A => \nb_send[3]_net_1\, B => \nb_send[4]_net_1\, 
        Y => \DWACT_FINC_E[1]\);
    
    un1_address_m49 : AX1C
      port map(A => \addr_data_vector[98]\, B => 
        \un1_state_12[4]\, C => \addr_data_vector[99]\, Y => 
        N_50_i_0);
    
    \address[9]\ : DFN1C0
      port map(D => \address_7[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[105]\);
    
    \address_RNO[18]\ : MX2
      port map(A => N_57_0, B => addr_data_f3(18), S => 
        \state_0[0]_net_1\, Y => \address_7[18]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \address_RNO[7]\ : MX2
      port map(A => N_1_i_0, B => addr_data_f3(7), S => 
        \state_0[0]_net_1\, Y => \address_7[7]\);
    
    un1_address_m48 : AX1C
      port map(A => \addr_data_vector[126]\, B => N_47, C => 
        \addr_data_vector[127]\, Y => N_49_i_0);
    
    \address[6]\ : DFN1C0
      port map(D => \address_7[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[102]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_59\ : OR2A
      port map(A => I_13_19, B => nb_burst_available(3), Y => 
        \ACT_LT4_E[8]\);
    
    \address_RNISVMA[4]\ : MX2C
      port map(A => addr_data_vector_0, B => 
        \addr_data_vector[100]\, S => sel_data_0(1), Y => N_1301);
    
    \FSM_SELECT_ADDRESS.state7_0_I_1\ : XNOR2
      port map(A => I_56_3, B => nb_burst_available(10), Y => 
        \DWACT_BL_EQUAL_0_E[4]\);
    
    status_full_err_RNO : AO1
      port map(A => \state[2]_net_1\, B => N_129, C => 
        un1_state_5_i_0, Y => N_110);
    
    \state_0[0]\ : DFN1C0
      port map(D => \state_RNIKABE[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state_0[0]_net_1\);
    
    \address_RNO[8]\ : MX2
      port map(A => N_15_0_i_0, B => addr_data_f3(8), S => 
        \state_0[0]_net_1\, Y => \address_7[8]\);
    
    \state_RNIQBSU8[3]\ : NOR3B
      port map(A => \state[3]_net_1\, B => state7, C => 
        un3_update_r, Y => address_0_sqmuxa);
    
    un1_address_m36 : NOR2A
      port map(A => \addr_data_vector[117]\, B => N_36_0, Y => 
        N_37_0);
    
    \state_RNI1KCD[1]\ : NOR2
      port map(A => \state[2]_net_1\, B => \state[1]_net_1\, Y
         => N_131);
    
    \address_RNIP245[28]\ : MX2C
      port map(A => addr_data_vector_24, B => 
        \addr_data_vector[124]\, S => sel_data(1), Y => N_911);
    
    un2_nb_send_next_I_52 : XOR2
      port map(A => N_7, B => \nb_send[9]_net_1\, Y => I_52_3);
    
    \address[11]\ : DFN1C0
      port map(D => \address_7[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[107]\);
    
    \address[31]\ : DFN1C0
      port map(D => \address_7[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[127]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_55\ : OR2A
      port map(A => nb_burst_available(2), B => I_9_19, Y => 
        \ACT_LT4_E[4]\);
    
    un1_address_m56 : AX1
      port map(A => N_29_0, B => \addr_data_vector[113]\, C => 
        \addr_data_vector[114]\, Y => N_57_0);
    
    \address_RNIE894[14]\ : MX2C
      port map(A => addr_data_vector_10, B => 
        \addr_data_vector[110]\, S => sel_data_0(1), Y => N_1283);
    
    \address_RNO[2]\ : MX2
      port map(A => N_40_i_0, B => addr_data_f3(2), S => 
        \state_0[0]_net_1\, Y => \address_7[2]\);
    
    \address_RNO[4]\ : MX2
      port map(A => N_51_i_0, B => addr_data_f3(4), S => 
        \state_0[0]_net_1\, Y => \address_7[4]\);
    
    un2_nb_send_next_I_19 : NOR2B
      port map(A => \nb_send[3]_net_1\, B => \DWACT_FINC_E[0]\, Y
         => N_30);
    
    \address_RNO[25]\ : MX2
      port map(A => N_61_0, B => addr_data_f3(25), S => 
        \state[0]_net_1\, Y => \address_7[25]\);
    
    \address[21]\ : DFN1C0
      port map(D => \address_7[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[117]\);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    un1_address_m62 : XNOR2
      port map(A => N_44, B => \addr_data_vector[123]\, Y => 
        N_63_0);
    
    un1_address_m32 : XNOR2
      port map(A => N_32_0, B => \addr_data_vector[115]\, Y => 
        N_33_0);
    
    un1_address_m12_e : OR3C
      port map(A => \addr_data_vector[100]\, B => N_69, C => 
        \addr_data_vector[101]\, Y => N_5_0);
    
    un2_nb_send_next_I_9 : XOR2
      port map(A => N_38, B => \nb_send[2]_net_1\, Y => I_9_19);
    
    \state[1]\ : DFN1C0
      port map(D => \state_RNO[1]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[1]_net_1\);
    
    un1_address_m24_m5_0_a2 : OR3C
      port map(A => m24_m5_0_a2_5, B => m24_m5_0_a2_4, C => 
        N_13_0, Y => N_25_0_i_0);
    
    \address[17]\ : DFN1C0
      port map(D => \address_7[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[113]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_52\ : OR2A
      port map(A => nb_burst_available(1), B => I_5_19, Y => 
        \ACT_LT4_E[1]\);
    
    un1_address_m65 : XOR2
      port map(A => N_47, B => \addr_data_vector[126]\, Y => 
        N_66_0);
    
    un1_address_m35 : OR3B
      port map(A => \addr_data_vector[115]\, B => 
        \addr_data_vector[116]\, C => N_32_0, Y => N_36_0);
    
    un1_address_m52 : XOR2
      port map(A => N_13_0, B => \addr_data_vector[103]\, Y => 
        N_1_i_0);
    
    un1_address_m24_m5_0_a2_5 : NOR3C
      port map(A => \addr_data_vector[107]\, B => 
        \addr_data_vector[106]\, C => m24_m5_0_a2_3, Y => 
        m24_m5_0_a2_5);
    
    \address_RNIM894[18]\ : MX2C
      port map(A => addr_data_vector_14, B => 
        \addr_data_vector[114]\, S => sel_data_0(1), Y => N_1287);
    
    un1_address_m24_m5_0_a2_3 : NOR2B
      port map(A => \addr_data_vector[108]\, B => 
        \addr_data_vector[109]\, Y => m24_m5_0_a2_3);
    
    \address[27]\ : DFN1C0
      port map(D => \address_7[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \addr_data_vector[123]\);
    
    \state_RNO[3]\ : NOR2A
      port map(A => \state[4]_net_1\, B => N_129, Y => 
        \state_RNO_0[3]\);
    
    un1_address_m21 : AX1C
      port map(A => \addr_data_vector[107]\, B => N_19_0, C => 
        \addr_data_vector[108]\, Y => N_22_0_i_0);
    
    \nb_send_RNO[4]\ : NOR2B
      port map(A => I_20_11, B => state7, Y => \nb_send_5[4]\);
    
    \nb_send_RNO[10]\ : NOR2B
      port map(A => I_56_3, B => state7, Y => \nb_send_5[10]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_18\ : OR2A
      port map(A => I_45_3, B => nb_burst_available(8), Y => N_29);
    
    un1_address_m55 : AX1C
      port map(A => \addr_data_vector[109]\, B => N_23_0, C => 
        \addr_data_vector[110]\, Y => N_56_0_i_0);
    
    \address_RNO[31]\ : MX2
      port map(A => N_49_i_0, B => addr_data_f3(31), S => 
        \state[0]_net_1\, Y => \address_7[31]\);
    
    \address_RNI2ONA[7]\ : MX2C
      port map(A => addr_data_vector_3, B => 
        \addr_data_vector[103]\, S => sel_data_0(1), Y => N_1290);
    
    \FSM_SELECT_ADDRESS.state7_0_I_61\ : AOI1A
      port map(A => \ACT_LT4_E[3]\, B => \ACT_LT4_E[6]\, C => 
        \ACT_LT4_E[10]\, Y => \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\);
    
    un1_address_m10_e : NOR3C
      port map(A => \addr_data_vector[98]\, B => 
        \un1_state_12[4]\, C => \addr_data_vector[99]\, Y => N_69);
    
    \FSM_SELECT_ADDRESS.state7_0_I_34\ : XNOR2
      port map(A => I_20_11, B => nb_burst_available(4), Y => 
        \DWACT_BL_EQUAL_0_E[0]\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_6\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E_0[0]\, B => 
        \DWACT_BL_EQUAL_0_E_0[1]\, C => \DWACT_BL_EQUAL_0_E[2]\, 
        Y => \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0]\);
    
    \address_RNO[12]\ : MX2
      port map(A => N_22_0_i_0, B => addr_data_f3(12), S => 
        \state_0[0]_net_1\, Y => \address_7[12]\);
    
    \update_r_RNI5KV4_0[0]\ : OR2
      port map(A => \update_r_i[0]\, B => \update_r[1]_net_1\, Y
         => \un1_state_12_3_0[4]\);
    
    un2_nb_send_next_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \nb_send[6]_net_1\, Y => N_17);
    
    un2_nb_send_next_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_12);
    
    \FSM_SELECT_ADDRESS.state7_0_I_3\ : XNOR2
      port map(A => I_45_3, B => nb_burst_available(8), Y => 
        \DWACT_BL_EQUAL_0_E[2]\);
    
    status_full_RNO : AO1A
      port map(A => state7, B => \state[3]_net_1\, C => 
        \state[2]_net_1\, Y => un1_state_11);
    
    \address_RNIHA45[31]\ : MX2C
      port map(A => addr_data_vector_27, B => 
        \addr_data_vector[127]\, S => sel_data(1), Y => N_914);
    
    \address[1]\ : DFN1E1C0
      port map(D => addr_data_f3(1), CLK => HCLK_c, CLR => 
        HRESETn_c, E => \state[0]_net_1\, Q => 
        addr_data_vector_61);
    
    \status_full\ : DFN1E1C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_11, Q => status_full(3));
    
    un1_address_m63 : AX1
      port map(A => N_44, B => \addr_data_vector[123]\, C => 
        \addr_data_vector[124]\, Y => N_64_0);
    
    un2_nb_send_next_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    \address_RNO[20]\ : MX2
      port map(A => N_35_0, B => addr_data_f3(20), S => 
        \state[0]_net_1\, Y => \address_7[20]\);
    
    un1_address_m46 : NOR2A
      port map(A => \addr_data_vector[125]\, B => N_46, Y => N_47);
    
    \nb_send[8]\ : DFN1E0C0
      port map(D => \nb_send_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[8]_net_1\);
    
    un1_address_m53 : AX1C
      port map(A => \addr_data_vector[105]\, B => N_16_0, C => 
        \addr_data_vector[106]\, Y => N_54_0_i_0);
    
    un1_address_m40_m6_0_a2_1 : NOR2B
      port map(A => \addr_data_vector[112]\, B => 
        \addr_data_vector[113]\, Y => m40_m6_0_a2_1);
    
    un1_address_m24_m5_0_a2_4 : NOR3C
      port map(A => \addr_data_vector[103]\, B => 
        \addr_data_vector[110]\, C => m24_m5_0_a2_1, Y => 
        m24_m5_0_a2_4);
    
    \nb_send[1]\ : DFN1E0C0
      port map(D => \nb_send_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_9, Q => \nb_send[1]_net_1\);
    
    \FSM_SELECT_ADDRESS.state7_0_I_60\ : AOI1A
      port map(A => \ACT_LT4_E[7]\, B => \ACT_LT4_E[8]\, C => 
        \ACT_LT4_E[5]\, Y => \ACT_LT4_E[10]\);
    
    \state_RNO_1[4]\ : OR3A
      port map(A => \state_0[0]_net_1\, B => \state[3]_net_1\, C
         => \state[2]_net_1\, Y => N_124);
    
    \address_RNO[15]\ : MX2
      port map(A => N_26_0_i_0, B => addr_data_f3(15), S => 
        \state_0[0]_net_1\, Y => \address_7[15]\);
    
    un2_nb_send_next_I_20 : XOR2
      port map(A => N_30, B => \nb_send[4]_net_1\, Y => I_20_11);
    
    \FSM_SELECT_ADDRESS.state7_0_I_68\ : AO1
      port map(A => \DWACT_CMPLE_PO2_DWACT_COMP0_E[1]\, B => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2]\, C => 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0]\, Y => 
        \DWACT_COMP0_E[2]\);
    
    un2_nb_send_next_I_16 : AND3
      port map(A => \nb_send[0]_net_1\, B => \nb_send[1]_net_1\, 
        C => \nb_send[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DMA2AHB is

    port( hburst_c           : out   std_logic_vector(2 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          un7_dmain          : in    std_logic_vector(66 to 66);
          hsize_c            : out   std_logic_vector(1 downto 0);
          AHB_Master_In_c_5  : in    std_logic;
          AHB_Master_In_c_4  : in    std_logic;
          AHB_Master_In_c_0  : in    std_logic;
          AHB_Master_In_c_3  : in    std_logic;
          haddr_c            : out   std_logic_vector(31 downto 0);
          hwrite_c           : out   std_logic;
          Ready              : out   std_logic;
          N_1012             : in    std_logic;
          Grant              : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          OKAY               : out   std_logic;
          Fault              : out   std_logic;
          N_1011             : in    std_logic;
          N_1013             : in    std_logic;
          N_43               : out   std_logic;
          time_select_0      : in    std_logic;
          N_960              : in    std_logic;
          N_959              : in    std_logic;
          N_958              : in    std_logic;
          N_957              : in    std_logic;
          N_964              : in    std_logic;
          N_963              : in    std_logic;
          N_962              : in    std_logic;
          N_961              : in    std_logic;
          N_955              : in    std_logic;
          N_954              : in    std_logic;
          N_953              : in    std_logic;
          N_952              : in    std_logic;
          N_951              : in    std_logic;
          N_950              : in    std_logic;
          N_949              : in    std_logic;
          N_948              : in    std_logic;
          N_947              : in    std_logic;
          N_956              : in    std_logic;
          N_965              : in    std_logic;
          N_966              : in    std_logic;
          N_967              : in    std_logic;
          N_968              : in    std_logic;
          N_969              : in    std_logic;
          N_970              : in    std_logic;
          N_971              : in    std_logic;
          N_972              : in    std_logic;
          N_973              : in    std_logic;
          N_974              : in    std_logic;
          N_975              : in    std_logic;
          N_976              : in    std_logic;
          N_977              : in    std_logic;
          HRESETn_c          : in    std_logic;
          N_978              : in    std_logic;
          HCLK_c             : in    std_logic
        );

end DMA2AHB;

architecture DEF_ARCH of DMA2AHB is 

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \htrans_12_i_o2_2_5[0]\, \htrans_12_i_o2_2_2[0]\, 
        \htrans_12_i_o2_2_4[0]\, \htrans_12_i_o2_2_0[0]\, N_183, 
        N_556_i_0, N_58_0, \Address_0_i_1[29]\, N_181, 
        \un1_AddressSave_0_sqmuxa_1_i_i[29]\, \Address_0_i_1[28]\, 
        N_179, N_37, \Address_0_i_1[26]\, N_177, N_35, 
        \Address_0_i_1[25]\, N_175, N_33_0, \Address_0_i_1[24]\, 
        N_173, N_55_0, \Address_0_i_1[23]\, N_128, N_556_i, 
        N_56_0, \Address_0_i_1[27]\, N_30, 
        \un1_AddressSave_0_sqmuxa_1_i_i[32]\, \Address_0_i_1[31]\, 
        N_28, N_42, \Address_0_i_1[30]\, N_13_0, N_580, N_15_0, 
        N_18_0, N_22_0, N_26_0, N_29_0, N_32_0, \haddr_c[24]\, 
        N_36, \haddr_c[25]\, N_39, \haddr_c[26]\, N_41, 
        \haddr_c[22]\, \haddr_c[23]\, \haddr_c[27]\, 
        \haddr_c[28]\, \haddr_c[29]\, \haddr_c[30]\, N_566, 
        \AddressPhase\, \AddressPhase_0\, N_191, hsize_0_sqmuxa_0, 
        N_756, N_754_0, \ReDataPhase\, N_553, N_753_0, N_555, 
        N_557, \Address_0_i_0[31]\, \AddressSave[31]_net_1\, 
        \Address_0_i_0[30]\, \AddressSave[30]_net_1\, 
        \Address_0_i_0[29]\, \AddressSave[29]_net_1\, 
        \Address_0_i_0[28]\, \AddressSave[28]_net_1\, 
        \Address_0_i_0[27]\, \AddressSave[27]_net_1\, 
        \Address_0_i_0[26]\, \AddressSave[26]_net_1\, 
        \Address_0_i_0[25]\, \AddressSave[25]_net_1\, 
        \Address_0_i_0[24]\, \AddressSave[24]_net_1\, 
        \Address_0_i_0[23]\, \AddressSave[23]_net_1\, 
        \Address_0_i_1[22]\, \Address_0_i_0[22]\, 
        \AddressSave[22]_net_1\, \Address_0_i_1[21]\, 
        \Address_0_i_0[21]\, \AddressSave[21]_net_1\, 
        \Address_0_i_1[20]\, \Address_0_i_0[20]\, 
        \AddressSave[20]_net_1\, \Address_0_i_1[19]\, 
        \Address_0_i_0[19]\, \AddressSave[19]_net_1\, 
        \Address_0_i_1[18]\, \Address_0_i_0[18]\, 
        \AddressSave[18]_net_1\, \Address_0_i_1[9]\, 
        \Address_0_i_0[9]\, \AddressSave[9]_net_1\, 
        \Address_0_i_1[0]\, \Address_0_i_0[0]\, 
        \AddressSave[0]_net_1\, \Address_0_i_1[1]\, N_753, 
        \Address_0_i_0[1]\, \AddressSave[1]_net_1\, N_754, 
        \Address_0_i_1[2]\, \Address_0_i_0[2]\, 
        \AddressSave[2]_net_1\, \Address_0_i_1[3]\, 
        \Address_0_i_0[3]\, \AddressSave[3]_net_1\, 
        \Address_0_i_1[4]\, \Address_0_i_0[4]\, 
        \AddressSave[4]_net_1\, \Address_0_i_1[5]\, 
        \Address_0_i_0[5]\, \AddressSave[5]_net_1\, 
        \Address_0_i_1[6]\, \Address_0_i_0[6]\, 
        \AddressSave[6]_net_1\, \Address_0_i_1[7]\, 
        \Address_0_i_0[7]\, \AddressSave[7]_net_1\, 
        \Address_0_i_1[8]\, \Address_0_i_0[8]\, 
        \AddressSave[8]_net_1\, \Address_0_i_1[14]\, 
        \Address_0_i_0[14]\, \AddressSave[14]_net_1\, 
        \Address_0_i_1[15]\, \Address_0_i_0[15]\, 
        \AddressSave[15]_net_1\, \Address_0_i_1[16]\, 
        \Address_0_i_0[16]\, \AddressSave[16]_net_1\, 
        \Address_0_i_1[17]\, \Address_0_i_0[17]\, 
        \AddressSave[17]_net_1\, \Address_0_i_1[10]\, 
        \Address_0_i_0[10]\, \AddressSave[10]_net_1\, 
        \Address_0_i_1[11]\, \Address_0_i_0[11]\, 
        \AddressSave[11]_net_1\, \Address_0_i_1[12]\, 
        \Address_0_i_0[12]\, \AddressSave[12]_net_1\, 
        \Address_0_i_1[13]\, \Address_0_i_0[13]\, 
        \AddressSave[13]_net_1\, \hsize_1_i_0[0]\, 
        BoundaryPhase_2_i_1, N_686, N_684, \hsize_1_i_0[1]\, 
        \htrans_12_i_2[0]\, \htrans_12_i_0[0]\, N_678, N_675, 
        \hsize_1_i_a5_0[1]\, \hsize_c[1]\, un1_ahbin_3_0_0, N_561, 
        \hburst_11_i_a2_i_a5_1[1]\, \ReAddrPhase\, 
        \hburst_11_0_a2_i_2[0]\, \hburst_11_0_a2_i_0[0]\, N_643, 
        N_563, \SingleAcc\, N_559, \un1_dmain_20_i_0\, 
        ActivePhase_1_sqmuxa_i_a5_0, \DataPhase\, DataPhase_2_i_0, 
        N_576, Fault_0_a5_0, \Address_RNO[13]_net_1\, 
        \un1_AddressSave_0_sqmuxa_1_i_i[14]\, 
        \Address_RNO[12]_net_1\, 
        \un1_AddressSave_0_sqmuxa_1_i_i[13]\, 
        \Address_RNO[11]_net_1\, 
        \un1_AddressSave_0_sqmuxa_1_i_i[12]\, 
        \Address_RNO[10]_net_1\, 
        \un1_AddressSave_0_sqmuxa_1_i_i[11]\, N_171, 
        \un1_AddressSave_0_sqmuxa_1_i_i[23]\, N_169, 
        \un1_AddressSave_0_sqmuxa_1_i_i[22]\, N_167, 
        \un1_AddressSave_0_sqmuxa_1_i_i[21]\, N_165, 
        \un1_AddressSave_0_sqmuxa_1_i_i[20]\, N_163, 
        \un1_AddressSave_0_sqmuxa_1_i_i[19]\, N_161, 
        \un1_AddressSave_0_sqmuxa_1_i_i[18]\, N_159, 
        \un1_AddressSave_0_sqmuxa_1_i_i[17]\, N_157, 
        \un1_AddressSave_0_sqmuxa_1_i_i[16]\, N_155, 
        \un1_AddressSave_0_sqmuxa_1_i_i[15]\, N_153, 
        \un1_AddressSave_0_sqmuxa_1_i_i[9]\, N_151, N_569, N_126, 
        \un1_AddressSave_0_sqmuxa_1_i_i[8]\, N_124, 
        \un1_AddressSave_0_sqmuxa_1_i_i[7]\, N_122, 
        \un1_AddressSave_0_sqmuxa_1_i_i[6]\, N_120, 
        \un1_AddressSave_0_sqmuxa_1_i_i[5]\, N_118, 
        \un1_AddressSave_0_sqmuxa_1_i_i[4]\, N_116, 
        \un1_AddressSave_0_sqmuxa_1_i_i[3]\, N_114, N_112, N_26, 
        \un1_AddressSave_0_sqmuxa_1_i_i[10]\, N_137_i_0, 
        \htrans_RNO_1[0]\, N_676, N_20, hwrite_2_sqmuxa, N_560, 
        hwrite_2_sqmuxa_1, N_758, N_149, N_147_i_0, 
        \BoundaryPhase_RNO_1\, N_685, N_635, \IdlePhase\, N_829, 
        N_567, N_760, N_682, N_554, N_189, N_737, N_196, N_193, 
        N_614, N_738, N_139, N_680, N_679, un1_ahbin_3, N_568, 
        N_639, N_56_i_0, N_330, N_592, N_331, N_593, N_332, N_594, 
        N_333, N_595, N_334, N_586, N_335, N_587, N_336, N_588, 
        N_337, N_589, N_338, N_613, N_339, N_590, N_340, N_615, 
        N_341, N_616, N_342, N_617, N_343, N_618, N_344, N_596, 
        N_345, N_597, N_346, N_598, hsize_0_sqmuxa, N_347, N_599, 
        N_348, N_600, N_349, N_601, N_350, N_602, N_351, N_603, 
        N_352, N_604, N_353, N_605, N_354, N_606, N_355, N_607, 
        N_356, N_608, N_357, N_609, N_358, N_610, N_359, N_611, 
        N_360, N_612, N_361, N_591, \haddr_c[2]\, N_5_0, 
        \haddr_c[3]\, \haddr_c[4]\, N_3_0, N_7_0, \haddr_c[5]\, 
        \haddr_c[6]\, N_9_0, \haddr_c[7]\, \haddr_c[8]\, 
        \haddr_c[10]\, \haddr_c[14]\, \haddr_c[16]\, 
        \haddr_c[17]\, \haddr_c[18]\, \haddr_c[19]\, 
        \haddr_c[20]\, \haddr_c[21]\, \haddr_c[9]\, \haddr_c[11]\, 
        \haddr_c[12]\, \haddr_c[13]\, \haddr_c[15]\, N_213, N_215, 
        N_217, N_219, N_221, N_225, N_259, N_261, N_263, N_279, 
        N_281, N_283, N_285, N_287, N_289, N_291, N_293, N_295, 
        \AddressSave_RNO[2]_net_1\, \AddressSave_RNO[3]_net_1\, 
        N_512, N_514, N_516, N_518, N_520, N_522, N_524, N_526, 
        N_528, N_530, N_532, N_534, \haddr_c[31]\, \haddr_c[0]\, 
        \haddr_c[1]\, \EarlyPhase\, N_562, N_325, N_53, N_48, 
        \BoundaryPhase\, Retry, N_761, N_102, SingleAcc_2_sqmuxa, 
        N_104, N_322, N_326, N_329, N_22, N_100, N_558, 
        \ActivePhase\, \WriteAcc\, N_582, N_130, N_24, N_327, 
        N_108, N_320, N_106, N_321, \hsize_c[0]\, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 

    hsize_c(1) <= \hsize_c[1]\;
    hsize_c(0) <= \hsize_c[0]\;
    haddr_c(31) <= \haddr_c[31]\;
    haddr_c(30) <= \haddr_c[30]\;
    haddr_c(29) <= \haddr_c[29]\;
    haddr_c(28) <= \haddr_c[28]\;
    haddr_c(27) <= \haddr_c[27]\;
    haddr_c(26) <= \haddr_c[26]\;
    haddr_c(25) <= \haddr_c[25]\;
    haddr_c(24) <= \haddr_c[24]\;
    haddr_c(23) <= \haddr_c[23]\;
    haddr_c(22) <= \haddr_c[22]\;
    haddr_c(21) <= \haddr_c[21]\;
    haddr_c(20) <= \haddr_c[20]\;
    haddr_c(19) <= \haddr_c[19]\;
    haddr_c(18) <= \haddr_c[18]\;
    haddr_c(17) <= \haddr_c[17]\;
    haddr_c(16) <= \haddr_c[16]\;
    haddr_c(15) <= \haddr_c[15]\;
    haddr_c(14) <= \haddr_c[14]\;
    haddr_c(13) <= \haddr_c[13]\;
    haddr_c(12) <= \haddr_c[12]\;
    haddr_c(11) <= \haddr_c[11]\;
    haddr_c(10) <= \haddr_c[10]\;
    haddr_c(9) <= \haddr_c[9]\;
    haddr_c(8) <= \haddr_c[8]\;
    haddr_c(7) <= \haddr_c[7]\;
    haddr_c(6) <= \haddr_c[6]\;
    haddr_c(5) <= \haddr_c[5]\;
    haddr_c(4) <= \haddr_c[4]\;
    haddr_c(3) <= \haddr_c[3]\;
    haddr_c(2) <= \haddr_c[2]\;
    haddr_c(1) <= \haddr_c[1]\;
    haddr_c(0) <= \haddr_c[0]\;

    \AHBOut.hwrite_RNO_0\ : OR2
      port map(A => \WriteAcc\, B => N_561, Y => N_680);
    
    \Address[16]\ : DFN1
      port map(D => N_159, CLK => HCLK_c, Q => \haddr_c[16]\);
    
    \Address[10]\ : DFN1
      port map(D => \Address_RNO[10]_net_1\, CLK => HCLK_c, Q => 
        \haddr_c[10]\);
    
    \Address_RNO_1[3]\ : OAI1
      port map(A => \AddressSave[3]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[3]\);
    
    \Address[30]\ : DFN1
      port map(D => N_28, CLK => HCLK_c, Q => \haddr_c[30]\);
    
    \AddressSave_RNO_0[30]\ : MX2
      port map(A => \AddressSave[30]_net_1\, B => N_612, S => 
        hsize_0_sqmuxa, Y => N_360);
    
    \AddressSave[8]\ : DFN1
      port map(D => N_283, CLK => HCLK_c, Q => 
        \AddressSave[8]_net_1\);
    
    \Address_RNO_1[0]\ : OAI1
      port map(A => \AddressSave[0]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[0]\);
    
    ReAddrPhase_RNIEV7K1 : NOR3B
      port map(A => N_829, B => \hburst_11_i_a2_i_a5_1[1]\, C => 
        N_554, Y => N_682);
    
    \DMAOut.Fault_0_a5_0\ : NOR2A
      port map(A => AHB_Master_In_c_4, B => AHB_Master_In_c_5, Y
         => Fault_0_a5_0);
    
    \AHBOut.hsize_RNO[1]\ : OA1B
      port map(A => N_569, B => \hsize_1_i_a5_0[1]\, C => 
        \hsize_1_i_0[1]\, Y => N_151);
    
    \Address_RNO[26]\ : OA1B
      port map(A => N_556_i_0, B => N_37, C => 
        \Address_0_i_1[26]\, Y => N_179);
    
    \AddressSave_RNO_0[12]\ : MX2
      port map(A => \AddressSave[12]_net_1\, B => N_617, S => 
        hsize_0_sqmuxa_0, Y => N_342);
    
    \AddressSave_RNO_1[1]\ : MX2
      port map(A => N_948, B => \haddr_c[1]\, S => 
        \AddressPhase_0\, Y => N_593);
    
    un1_AddressSave_0_sqmuxa_1_m55 : AX1C
      port map(A => \haddr_c[26]\, B => N_36, C => \haddr_c[27]\, 
        Y => N_56_0);
    
    EarlyPhase_RNIP1701 : NOR3B
      port map(A => N_561, B => AHB_Master_In_c_3, C => N_1011, Y
         => N_738);
    
    \Address_RNO[1]\ : OA1B
      port map(A => \haddr_c[1]\, B => N_556_i, C => 
        \Address_0_i_1[1]\, Y => N_114);
    
    \AddressSave_RNO_0[10]\ : MX2
      port map(A => \AddressSave[10]_net_1\, B => N_615, S => 
        hsize_0_sqmuxa_0, Y => N_340);
    
    \AddressSave_RNO_0[27]\ : MX2
      port map(A => \AddressSave[27]_net_1\, B => N_609, S => 
        hsize_0_sqmuxa, Y => N_357);
    
    \AddressSave[15]\ : DFN1
      port map(D => N_287, CLK => HCLK_c, Q => 
        \AddressSave[15]_net_1\);
    
    un1_AddressSave_0_sqmuxa_1_m50 : XOR2
      port map(A => N_13_0, B => \haddr_c[12]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[13]\);
    
    \Address[26]\ : DFN1
      port map(D => N_179, CLK => HCLK_c, Q => \haddr_c[26]\);
    
    \Address[20]\ : DFN1
      port map(D => N_167, CLK => HCLK_c, Q => \haddr_c[20]\);
    
    \AddressSave[12]\ : DFN1
      port map(D => N_285, CLK => HCLK_c, Q => 
        \AddressSave[12]_net_1\);
    
    \AddressSave_RNO_1[16]\ : MX2
      port map(A => N_963, B => \haddr_c[16]\, S => 
        \AddressPhase_0\, Y => N_598);
    
    \Address_RNO_1[8]\ : OAI1
      port map(A => \AddressSave[8]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[8]\);
    
    BoundaryPhase_RNO : NOR3C
      port map(A => BoundaryPhase_2_i_1, B => 
        \BoundaryPhase_RNO_1\, C => N_685, Y => N_147_i_0);
    
    un1_AddressSave_0_sqmuxa_1_m31 : NOR3C
      port map(A => \haddr_c[22]\, B => N_29_0, C => 
        \haddr_c[23]\, Y => N_32_0);
    
    IdlePhase_RNO : NOR2B
      port map(A => N_326, B => HRESETn_c, Y => N_100);
    
    un1_AddressSave_0_sqmuxa_1_m47 : XNOR2
      port map(A => N_9_0, B => \haddr_c[9]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[10]\);
    
    \AHBOut.hsize[1]\ : DFN1
      port map(D => N_151, CLK => HCLK_c, Q => \hsize_c[1]\);
    
    ActivePhase_RNO_2 : OR2
      port map(A => \DataPhase\, B => \AddressPhase_0\, Y => 
        ActivePhase_1_sqmuxa_i_a5_0);
    
    \AHBOut.hburst_RNO_1[0]\ : AOI1B
      port map(A => \SingleAcc\, B => N_559, C => 
        AHB_Master_In_c_0, Y => \hburst_11_0_a2_i_0[0]\);
    
    \Address_RNO_0[11]\ : AO1D
      port map(A => N_958, B => N_753, C => \Address_0_i_0[11]\, 
        Y => \Address_0_i_1[11]\);
    
    \Address_RNO_0[8]\ : AO1D
      port map(A => N_955, B => N_753, C => \Address_0_i_0[8]\, Y
         => \Address_0_i_1[8]\);
    
    \Address_RNO_1[21]\ : OAI1
      port map(A => \AddressSave[21]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[21]\);
    
    \AHBOut.hwrite\ : DFN1E1
      port map(D => N_139, CLK => HCLK_c, E => N_130, Q => 
        hwrite_c);
    
    \Address[12]\ : DFN1
      port map(D => \Address_RNO[12]_net_1\, CLK => HCLK_c, Q => 
        \haddr_c[12]\);
    
    \AddressSave[23]\ : DFN1
      port map(D => N_526, CLK => HCLK_c, Q => 
        \AddressSave[23]_net_1\);
    
    \AddressSave_RNO_0[8]\ : MX2
      port map(A => \AddressSave[8]_net_1\, B => N_613, S => 
        hsize_0_sqmuxa_0, Y => N_338);
    
    \AddressSave_RNO_1[31]\ : MX2
      port map(A => N_978, B => \haddr_c[31]\, S => 
        \AddressPhase_0\, Y => N_591);
    
    \AddressSave_RNO[5]\ : NOR2B
      port map(A => N_335, B => HRESETn_c, Y => N_281);
    
    \Address_RNO_1[11]\ : OAI1
      port map(A => \AddressSave[11]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[11]\);
    
    \AddressSave_RNO[18]\ : NOR2B
      port map(A => N_348, B => HRESETn_c, Y => N_524);
    
    un1_AddressSave_0_sqmuxa_1_m41 : XOR2
      port map(A => N_41, B => \haddr_c[30]\, Y => N_42);
    
    \Address_RNO[29]\ : OA1B
      port map(A => N_556_i_0, B => N_58_0, C => 
        \Address_0_i_1[29]\, Y => N_183);
    
    \AddressSave_RNO_1[28]\ : MX2A
      port map(A => N_975, B => \haddr_c[28]\, S => 
        \AddressPhase\, Y => N_610);
    
    WriteAcc_RNO : NOR2B
      port map(A => N_321, B => HRESETn_c, Y => N_106);
    
    \AddressSave_RNO[11]\ : NOR2B
      port map(A => N_341, B => HRESETn_c, Y => N_518);
    
    SingleAcc_RNO : NOR2B
      port map(A => N_322, B => HRESETn_c, Y => N_104);
    
    ReAddrPhase_RNO_1 : OA1B
      port map(A => \AddressPhase\, B => \ReAddrPhase\, C => 
        AHB_Master_In_c_3, Y => N_53);
    
    \Address[22]\ : DFN1
      port map(D => N_171, CLK => HCLK_c, Q => \haddr_c[22]\);
    
    \Address_RNO[23]\ : OA1B
      port map(A => N_556_i_0, B => N_55_0, C => 
        \Address_0_i_1[23]\, Y => N_173);
    
    \Address[2]\ : DFN1
      port map(D => N_116, CLK => HCLK_c, Q => \haddr_c[2]\);
    
    \Address_RNO_1[7]\ : OAI1
      port map(A => \AddressSave[7]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[7]\);
    
    \Address_RNO[24]\ : OA1B
      port map(A => N_556_i_0, B => N_33_0, C => 
        \Address_0_i_1[24]\, Y => N_175);
    
    \Address_RNO[10]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[11]\, C => 
        \Address_0_i_1[10]\, Y => \Address_RNO[10]_net_1\);
    
    \AddressSave[20]\ : DFN1
      port map(D => N_225, CLK => HCLK_c, Q => 
        \AddressSave[20]_net_1\);
    
    \Address_RNO_1[30]\ : OAI1
      port map(A => \AddressSave[30]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[30]\);
    
    \AddressSave_RNO_1[3]\ : MX2
      port map(A => N_950, B => \haddr_c[3]\, S => 
        \AddressPhase_0\, Y => N_595);
    
    \AddressSave_RNO_1[19]\ : MX2
      port map(A => N_966, B => \haddr_c[19]\, S => 
        \AddressPhase_0\, Y => N_601);
    
    AddressPhase_RNI6S87 : OR2B
      port map(A => \AddressPhase\, B => AHB_Master_In_c_3, Y => 
        N_566);
    
    ActivePhase_RNIS2FG1 : AO1
      port map(A => N_582, B => AHB_Master_In_c_3, C => N_563, Y
         => N_130);
    
    EarlyPhase_RNO_1 : AO1C
      port map(A => AHB_Master_In_c_0, B => N_568, C => 
        un1_ahbin_3_0_0, Y => un1_ahbin_3);
    
    \AddressSave_RNO_1[24]\ : MX2
      port map(A => N_971, B => \haddr_c[24]\, S => 
        \AddressPhase\, Y => N_606);
    
    \DMAOut.Ready_RNO\ : NOR3C
      port map(A => HRESETn_c, B => AHB_Master_In_c_3, C => 
        \DataPhase\, Y => N_196);
    
    BoundaryPhase_RNO_2 : OR2A
      port map(A => N_555, B => N_553, Y => N_685);
    
    \AddressSave_RNO[25]\ : NOR2B
      port map(A => N_355, B => HRESETn_c, Y => N_530);
    
    \AddressSave_RNO_1[23]\ : MX2
      port map(A => N_970, B => \haddr_c[23]\, S => 
        \AddressPhase\, Y => N_605);
    
    \AHBOut.hbusreq_i_0_a2\ : NOR2A
      port map(A => un7_dmain(66), B => N_1011, Y => N_761);
    
    \Address_RNO[9]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[10]\, C => 
        \Address_0_i_1[9]\, Y => N_26);
    
    \Address[5]\ : DFN1
      port map(D => N_122, CLK => HCLK_c, Q => \haddr_c[5]\);
    
    \AddressSave[30]\ : DFN1
      port map(D => N_532, CLK => HCLK_c, Q => 
        \AddressSave[30]_net_1\);
    
    \Address[15]\ : DFN1
      port map(D => N_157, CLK => HCLK_c, Q => \haddr_c[15]\);
    
    \AHBOut.hburst[2]\ : DFN1E1
      port map(D => N_682, CLK => HCLK_c, E => N_130, Q => 
        hburst_c(2));
    
    \Address_RNO_0[9]\ : AO1D
      port map(A => N_956, B => N_753_0, C => \Address_0_i_0[9]\, 
        Y => \Address_0_i_1[9]\);
    
    \Address[13]\ : DFN1
      port map(D => \Address_RNO[13]_net_1\, CLK => HCLK_c, Q => 
        \haddr_c[13]\);
    
    \AddressSave_RNO_1[15]\ : MX2
      port map(A => N_962, B => \haddr_c[15]\, S => 
        \AddressPhase_0\, Y => N_597);
    
    \AddressSave_RNO_1[11]\ : MX2
      port map(A => N_958, B => \haddr_c[11]\, S => 
        \AddressPhase\, Y => N_616);
    
    \AddressSave_RNO_0[18]\ : MX2
      port map(A => \AddressSave[18]_net_1\, B => N_600, S => 
        hsize_0_sqmuxa, Y => N_348);
    
    \AddressSave[6]\ : DFN1
      port map(D => N_215, CLK => HCLK_c, Q => 
        \AddressSave[6]_net_1\);
    
    un1_AddressSave_0_sqmuxa_1_m24 : AX1C
      port map(A => \haddr_c[18]\, B => N_22_0, C => 
        \haddr_c[19]\, Y => \un1_AddressSave_0_sqmuxa_1_i_i[20]\);
    
    \AHBOut.hsize_RNO_1[1]\ : OR2
      port map(A => \hsize_c[1]\, B => \AddressPhase_0\, Y => 
        \hsize_1_i_a5_0[1]\);
    
    \Address_RNO_1[4]\ : OAI1
      port map(A => \AddressSave[4]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[4]\);
    
    ReDataPhase_RNIORDS : OA1B
      port map(A => N_555, B => \ReDataPhase\, C => N_553, Y => 
        N_556_i);
    
    \Address[19]\ : DFN1
      port map(D => N_165, CLK => HCLK_c, Q => \haddr_c[19]\);
    
    ActivePhase_RNII8GG : OR2A
      port map(A => N_1011, B => \ActivePhase\, Y => N_554);
    
    BoundaryPhase_RNO_0 : NOR3C
      port map(A => N_686, B => HRESETn_c, C => N_684, Y => 
        BoundaryPhase_2_i_1);
    
    \Address[25]\ : DFN1
      port map(D => N_177, CLK => HCLK_c, Q => \haddr_c[25]\);
    
    un1_AddressSave_0_sqmuxa_1_m12 : NOR3C
      port map(A => \haddr_c[10]\, B => N_580, C => \haddr_c[11]\, 
        Y => N_13_0);
    
    \Address_RNO_0[27]\ : AO1A
      port map(A => N_753_0, B => N_974, C => \Address_0_i_0[27]\, 
        Y => \Address_0_i_1[27]\);
    
    \AddressSave_RNO[7]\ : NOR2B
      port map(A => N_337, B => HRESETn_c, Y => N_217);
    
    ActivePhase_RNIHBAN : OR2
      port map(A => N_554, B => N_553, Y => N_756);
    
    \Address[23]\ : DFN1
      port map(D => N_173, CLK => HCLK_c, Q => \haddr_c[23]\);
    
    \AddressSave_RNO_1[7]\ : MX2
      port map(A => N_954, B => \haddr_c[7]\, S => 
        \AddressPhase_0\, Y => N_589);
    
    \AHBOut.htrans[1]\ : DFN1E1
      port map(D => N_193, CLK => HCLK_c, E => N_189, Q => 
        htrans_c(1));
    
    DataPhase_RNI0SGJ_0 : AO1C
      port map(A => N_760, B => N_558, C => HRESETn_c, Y => N_563);
    
    AddressPhase_RNIDRDU1 : NOR3
      port map(A => N_563, B => N_614, C => N_738, Y => N_191);
    
    WriteAcc_RNO_0 : MX2
      port map(A => \WriteAcc\, B => N_1012, S => hwrite_2_sqmuxa, 
        Y => N_321);
    
    \AddressSave_RNO[29]\ : NOR2B
      port map(A => N_359, B => HRESETn_c, Y => N_295);
    
    \AddressSave_RNO_0[14]\ : MX2
      port map(A => \AddressSave[14]_net_1\, B => N_596, S => 
        hsize_0_sqmuxa_0, Y => N_344);
    
    \Address[29]\ : DFN1
      port map(D => N_183, CLK => HCLK_c, Q => \haddr_c[29]\);
    
    \Address_RNIQTTQ[4]\ : NOR3C
      port map(A => \haddr_c[4]\, B => \haddr_c[3]\, C => 
        \htrans_12_i_o2_2_0[0]\, Y => \htrans_12_i_o2_2_4[0]\);
    
    \Address[18]\ : DFN1
      port map(D => N_163, CLK => HCLK_c, Q => \haddr_c[18]\);
    
    \AddressSave_RNO[10]\ : NOR2B
      port map(A => N_340, B => HRESETn_c, Y => N_516);
    
    \AddressSave[16]\ : DFN1
      port map(D => N_520, CLK => HCLK_c, Q => 
        \AddressSave[16]_net_1\);
    
    \AddressSave_RNO_1[26]\ : MX2A
      port map(A => N_973, B => \haddr_c[26]\, S => 
        \AddressPhase\, Y => N_608);
    
    \AddressSave_RNO_0[13]\ : MX2
      port map(A => \AddressSave[13]_net_1\, B => N_618, S => 
        hsize_0_sqmuxa_0, Y => N_343);
    
    ActivePhase_RNO : NOR2B
      port map(A => N_320, B => HRESETn_c, Y => N_108);
    
    \Address_RNO[21]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[22]\, C => 
        \Address_0_i_1[21]\, Y => N_169);
    
    \Address_RNO[16]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[17]\, C => 
        \Address_0_i_1[16]\, Y => N_159);
    
    SingleAcc_RNO_1 : NOR3C
      port map(A => AHB_Master_In_c_0, B => N_561, C => 
        un7_dmain(66), Y => SingleAcc_2_sqmuxa);
    
    \Address_RNO_0[30]\ : AO1D
      port map(A => N_977, B => N_753_0, C => \Address_0_i_0[30]\, 
        Y => \Address_0_i_1[30]\);
    
    \Address_RNO_0[24]\ : AO1D
      port map(A => N_971, B => N_753_0, C => \Address_0_i_0[24]\, 
        Y => \Address_0_i_1[24]\);
    
    un1_AddressSave_0_sqmuxa_1_m2 : OR2A
      port map(A => \haddr_c[2]\, B => N_566, Y => N_3_0);
    
    \Address_RNO_0[25]\ : AO1D
      port map(A => N_972, B => N_753_0, C => \Address_0_i_0[25]\, 
        Y => \Address_0_i_1[25]\);
    
    \Address[0]\ : DFN1
      port map(D => N_112, CLK => HCLK_c, Q => \haddr_c[0]\);
    
    ReDataPhase_RNIHO18 : OR2A
      port map(A => \ReDataPhase\, B => N_553, Y => N_754);
    
    \AddressSave_RNO[22]\ : NOR2B
      port map(A => N_352, B => HRESETn_c, Y => N_291);
    
    DataPhase_RNIFGQC : NOR2A
      port map(A => AHB_Master_In_c_5, B => N_760, Y => Retry);
    
    BoundaryPhase_RNO_1 : OR2
      port map(A => N_580, B => \BoundaryPhase\, Y => 
        \BoundaryPhase_RNO_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \AddressSave_RNO_0[6]\ : MX2
      port map(A => \AddressSave[6]_net_1\, B => N_588, S => 
        hsize_0_sqmuxa_0, Y => N_336);
    
    \AHBOut.hsize_RNO_2[1]\ : OAI1
      port map(A => AHB_Master_In_c_3, B => \hsize_c[1]\, C => 
        HRESETn_c, Y => \hsize_1_i_0[1]\);
    
    \AHBOut.hburst_RNO_0[0]\ : NOR3B
      port map(A => \hburst_11_0_a2_i_0[0]\, B => N_643, C => 
        N_563, Y => \hburst_11_0_a2_i_2[0]\);
    
    \AddressSave_RNO[16]\ : NOR2B
      port map(A => N_346, B => HRESETn_c, Y => N_520);
    
    \Address_RNO[27]\ : OA1B
      port map(A => N_556_i, B => N_56_0, C => 
        \Address_0_i_1[27]\, Y => N_128);
    
    \Address[4]\ : DFN1
      port map(D => N_120, CLK => HCLK_c, Q => \haddr_c[4]\);
    
    \Address[28]\ : DFN1
      port map(D => N_181, CLK => HCLK_c, Q => \haddr_c[28]\);
    
    \AHBOut.htrans_RNO_5[0]\ : OAI1
      port map(A => \ReAddrPhase\, B => N_1011, C => 
        \BoundaryPhase\, Y => N_675);
    
    \AddressSave_RNO[23]\ : NOR2B
      port map(A => N_353, B => HRESETn_c, Y => N_526);
    
    un1_AddressSave_0_sqmuxa_1_m49 : AX1C
      port map(A => \haddr_c[10]\, B => N_580, C => \haddr_c[11]\, 
        Y => \un1_AddressSave_0_sqmuxa_1_i_i[12]\);
    
    un1_AddressSave_0_sqmuxa_1_m35 : NOR3C
      port map(A => \haddr_c[24]\, B => N_32_0, C => 
        \haddr_c[25]\, Y => N_36);
    
    \Address_RNO_0[3]\ : AO1D
      port map(A => N_950, B => N_753, C => \Address_0_i_0[3]\, Y
         => \Address_0_i_1[3]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un1_AddressSave_0_sqmuxa_1_m52 : AX1C
      port map(A => \haddr_c[14]\, B => N_15_0, C => 
        \haddr_c[15]\, Y => \un1_AddressSave_0_sqmuxa_1_i_i[16]\);
    
    EarlyPhase : DFN1
      port map(D => N_24, CLK => HCLK_c, Q => \EarlyPhase\);
    
    \Address_RNO_1[31]\ : OAI1
      port map(A => \AddressSave[31]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[31]\);
    
    \AddressSave_RNO[4]\ : NOR2B
      port map(A => N_334, B => HRESETn_c, Y => N_512);
    
    un1_AddressSave_0_sqmuxa_1_m18 : XOR2
      port map(A => N_18_0, B => \haddr_c[16]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[17]\);
    
    \Address_RNO_0[4]\ : AO1D
      port map(A => N_951, B => N_753, C => \Address_0_i_0[4]\, Y
         => \Address_0_i_1[4]\);
    
    \Address_RNO_0[5]\ : AO1D
      port map(A => N_952, B => N_753, C => \Address_0_i_0[5]\, Y
         => \Address_0_i_1[5]\);
    
    \AHBOut.hsize[0]\ : DFN1
      port map(D => N_149, CLK => HCLK_c, Q => \hsize_c[0]\);
    
    \Address_RNO_0[17]\ : AO1D
      port map(A => N_964, B => N_753, C => \Address_0_i_0[17]\, 
        Y => \Address_0_i_1[17]\);
    
    \AddressSave_RNO_1[2]\ : MX2
      port map(A => N_949, B => \haddr_c[2]\, S => 
        \AddressPhase_0\, Y => N_594);
    
    ReAddrPhase_RNO : NOR2B
      port map(A => N_325, B => HRESETn_c, Y => N_102);
    
    \AddressSave_RNO_1[17]\ : MX2
      port map(A => N_964, B => \haddr_c[17]\, S => 
        \AddressPhase_0\, Y => N_599);
    
    \Address_RNO_1[27]\ : OAI1
      port map(A => \AddressSave[27]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[27]\);
    
    \AHBMaster.AHBOut.hwrite_8_iv_i_o5\ : OR2B
      port map(A => AHB_Master_In_c_3, B => AHB_Master_In_c_0, Y
         => N_553);
    
    un1_AddressSave_0_sqmuxa_1_m45 : AX1
      port map(A => N_5_0, B => \haddr_c[5]\, C => \haddr_c[6]\, 
        Y => \un1_AddressSave_0_sqmuxa_1_i_i[7]\);
    
    \Address_RNI2UUQ[8]\ : NOR3C
      port map(A => \haddr_c[8]\, B => \haddr_c[7]\, C => 
        \htrans_12_i_o2_2_2[0]\, Y => \htrans_12_i_o2_2_5[0]\);
    
    \Address_RNO[19]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[20]\, C => 
        \Address_0_i_1[19]\, Y => N_165);
    
    \AddressSave_RNO_0[16]\ : MX2
      port map(A => \AddressSave[16]_net_1\, B => N_598, S => 
        hsize_0_sqmuxa, Y => N_346);
    
    \Address_RNO_1[17]\ : OAI1
      port map(A => \AddressSave[17]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[17]\);
    
    \AHBOut.hburst[0]\ : DFN1E1
      port map(D => N_56_i_0, CLK => HCLK_c, E => N_130, Q => 
        hburst_c(0));
    
    \AddressSave[9]\ : DFN1
      port map(D => N_514, CLK => HCLK_c, Q => 
        \AddressSave[9]_net_1\);
    
    un1_AddressSave_0_sqmuxa_1_m40 : NOR3C
      port map(A => \haddr_c[28]\, B => N_39, C => \haddr_c[29]\, 
        Y => N_41);
    
    IdlePhase_0_sqmuxa_0_o2 : OR2
      port map(A => AHB_Master_In_c_5, B => AHB_Master_In_c_4, Y
         => N_558);
    
    \AddressSave_RNO_1[29]\ : MX2
      port map(A => N_976, B => \haddr_c[29]\, S => 
        \AddressPhase\, Y => N_611);
    
    \AddressSave_RNO[2]\ : NOR2B
      port map(A => N_332, B => HRESETn_c, Y => 
        \AddressSave_RNO[2]_net_1\);
    
    \Address_RNO[13]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[14]\, C => 
        \Address_0_i_1[13]\, Y => \Address_RNO[13]_net_1\);
    
    \Address_RNO_0[14]\ : AO1D
      port map(A => N_961, B => N_753, C => \Address_0_i_0[14]\, 
        Y => \Address_0_i_1[14]\);
    
    \Address[14]\ : DFN1
      port map(D => N_155, CLK => HCLK_c, Q => \haddr_c[14]\);
    
    \AddressSave[29]\ : DFN1
      port map(D => N_295, CLK => HCLK_c, Q => 
        \AddressSave[29]_net_1\);
    
    \Address_RNO_0[15]\ : AO1D
      port map(A => N_962, B => N_753, C => \Address_0_i_0[15]\, 
        Y => \Address_0_i_1[15]\);
    
    \Address_RNO_1[24]\ : OAI1
      port map(A => \AddressSave[24]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[24]\);
    
    \AddressSave_RNO_0[1]\ : MX2
      port map(A => \AddressSave[1]_net_1\, B => N_593, S => 
        hsize_0_sqmuxa_0, Y => N_331);
    
    \IdlePhase_RNI03G71\ : OA1C
      port map(A => N_761, B => N_559, C => \IdlePhase\, Y => 
        IdlePhase_RNI03G71);
    
    \Address_RNO_1[25]\ : OAI1
      port map(A => \AddressSave[25]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[25]\);
    
    \Address_RNO[14]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[15]\, C => 
        \Address_0_i_1[14]\, Y => N_155);
    
    \Address_RNO_1[14]\ : OAI1
      port map(A => \AddressSave[14]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[14]\);
    
    \Address_RNIV6FD[6]\ : NOR2B
      port map(A => \haddr_c[5]\, B => \haddr_c[6]\, Y => 
        \htrans_12_i_o2_2_2[0]\);
    
    DataPhase_RNIGGQC : OR2B
      port map(A => N_558, B => \DataPhase\, Y => N_737);
    
    \Address_RNO_1[15]\ : OAI1
      port map(A => \AddressSave[15]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[15]\);
    
    \AddressSave[11]\ : DFN1
      port map(D => N_518, CLK => HCLK_c, Q => 
        \AddressSave[11]_net_1\);
    
    \AddressSave_RNO_1[25]\ : MX2
      port map(A => N_972, B => \haddr_c[25]\, S => 
        \AddressPhase\, Y => N_607);
    
    \AddressSave_RNO_1[21]\ : MX2
      port map(A => N_968, B => \haddr_c[21]\, S => 
        \AddressPhase_0\, Y => N_603);
    
    \Address[24]\ : DFN1
      port map(D => N_175, CLK => HCLK_c, Q => \haddr_c[24]\);
    
    \Address_RNO_0[22]\ : AO1D
      port map(A => N_969, B => N_753_0, C => \Address_0_i_0[22]\, 
        Y => \Address_0_i_1[22]\);
    
    \AddressSave[1]\ : DFN1
      port map(D => N_279, CLK => HCLK_c, Q => 
        \AddressSave[1]_net_1\);
    
    \AHBOut.hwrite_RNO\ : NOR3C
      port map(A => N_193, B => N_680, C => N_679, Y => N_139);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Address_RNO_0[31]\ : AO1D
      port map(A => N_978, B => N_753_0, C => \Address_0_i_0[31]\, 
        Y => \Address_0_i_1[31]\);
    
    \AddressSave[25]\ : DFN1
      port map(D => N_530, CLK => HCLK_c, Q => 
        \AddressSave[25]_net_1\);
    
    un1_AddressSave_0_sqmuxa_1_m27 : AX1C
      port map(A => \haddr_c[20]\, B => N_26_0, C => 
        \haddr_c[21]\, Y => \un1_AddressSave_0_sqmuxa_1_i_i[22]\);
    
    \AddressSave[22]\ : DFN1
      port map(D => N_291, CLK => HCLK_c, Q => 
        \AddressSave[22]_net_1\);
    
    \AddressSave_RNO_0[19]\ : MX2
      port map(A => \AddressSave[19]_net_1\, B => N_601, S => 
        hsize_0_sqmuxa, Y => N_349);
    
    ReDataPhase_RNIORDS_0 : OA1B
      port map(A => N_555, B => \ReDataPhase\, C => N_553, Y => 
        N_556_i_0);
    
    \AddressSave_RNO_0[31]\ : MX2
      port map(A => \AddressSave[31]_net_1\, B => N_591, S => 
        hsize_0_sqmuxa, Y => N_361);
    
    \AddressSave_RNO[1]\ : NOR2B
      port map(A => N_331, B => HRESETn_c, Y => N_279);
    
    \Address[8]\ : DFN1
      port map(D => N_153, CLK => HCLK_c, Q => \haddr_c[8]\);
    
    \Address_RNO_0[1]\ : AO1D
      port map(A => N_948, B => N_753, C => \Address_0_i_0[1]\, Y
         => \Address_0_i_1[1]\);
    
    un1_AddressSave_0_sqmuxa_1_m21 : NOR3C
      port map(A => \haddr_c[16]\, B => N_18_0, C => 
        \haddr_c[17]\, Y => N_22_0);
    
    BoundaryPhase : DFN1
      port map(D => N_147_i_0, CLK => HCLK_c, Q => 
        \BoundaryPhase\);
    
    \AddressSave_RNO_0[7]\ : MX2
      port map(A => \AddressSave[7]_net_1\, B => N_589, S => 
        hsize_0_sqmuxa_0, Y => N_337);
    
    ReAddrPhase_RNO_2 : AO1A
      port map(A => N_557, B => \ReAddrPhase\, C => Retry, Y => 
        N_48);
    
    EarlyPhase_RNILB3D : NOR2
      port map(A => N_559, B => \EarlyPhase\, Y => N_561);
    
    \AddressSave_RNO[24]\ : NOR2B
      port map(A => N_354, B => HRESETn_c, Y => N_528);
    
    \AHBOut.htrans_RNO_0[0]\ : NOR3C
      port map(A => \htrans_12_i_0[0]\, B => N_678, C => N_675, Y
         => \htrans_12_i_2[0]\);
    
    \AddressSave_RNO_1[9]\ : MX2
      port map(A => N_956, B => \haddr_c[9]\, S => 
        \AddressPhase_0\, Y => N_590);
    
    \AHBOut.hburst_RNO_2[0]\ : OR2B
      port map(A => un7_dmain(66), B => N_561, Y => N_643);
    
    \Address_RNO[6]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[7]\, C => 
        \Address_0_i_1[6]\, Y => N_124);
    
    IdlePhase : DFN1
      port map(D => N_100, CLK => HCLK_c, Q => \IdlePhase\);
    
    \AddressSave_RNO_0[15]\ : MX2
      port map(A => \AddressSave[15]_net_1\, B => N_597, S => 
        hsize_0_sqmuxa_0, Y => N_345);
    
    \AddressSave_RNO_0[11]\ : MX2
      port map(A => \AddressSave[11]_net_1\, B => N_616, S => 
        hsize_0_sqmuxa_0, Y => N_341);
    
    ReAddrPhase : DFN1
      port map(D => N_102, CLK => HCLK_c, Q => \ReAddrPhase\);
    
    \Address_RNO[28]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[29]\, C => 
        \Address_0_i_1[28]\, Y => N_181);
    
    \Address_RNO[11]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[12]\, C => 
        \Address_0_i_1[11]\, Y => \Address_RNO[11]_net_1\);
    
    \Address_RNO_0[12]\ : AO1D
      port map(A => N_959, B => N_753, C => \Address_0_i_0[12]\, 
        Y => \Address_0_i_1[12]\);
    
    \AddressSave_RNO_1[5]\ : MX2
      port map(A => N_952, B => \haddr_c[5]\, S => 
        \AddressPhase_0\, Y => N_587);
    
    DataPhase_RNO_0 : OAI1
      port map(A => AHB_Master_In_c_3, B => N_576, C => HRESETn_c, 
        Y => DataPhase_2_i_0);
    
    \Address_RNO_1[22]\ : OAI1
      port map(A => \AddressSave[22]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[22]\);
    
    \Address_RNO[17]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[18]\, C => 
        \Address_0_i_1[17]\, Y => N_161);
    
    \AddressSave_RNO_0[0]\ : MX2
      port map(A => \AddressSave[0]_net_1\, B => N_592, S => 
        hsize_0_sqmuxa_0, Y => N_330);
    
    \AddressSave_RNO[31]\ : NOR2B
      port map(A => N_361, B => HRESETn_c, Y => N_534);
    
    IdlePhase_RNI9HPU : NOR3
      port map(A => N_635, B => \IdlePhase\, C => N_1013, Y => 
        N_43);
    
    \Address_RNO[5]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[6]\, C => 
        \Address_0_i_1[5]\, Y => N_122);
    
    \AddressSave[17]\ : DFN1
      port map(D => N_522, CLK => HCLK_c, Q => 
        \AddressSave[17]_net_1\);
    
    \Address_RNO_1[12]\ : OAI1
      port map(A => \AddressSave[12]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[12]\);
    
    \AddressSave_RNO_1[27]\ : MX2A
      port map(A => N_974, B => \haddr_c[27]\, S => 
        \AddressPhase\, Y => N_609);
    
    \AddressSave_RNO[15]\ : NOR2B
      port map(A => N_345, B => HRESETn_c, Y => N_287);
    
    \AddressSave[4]\ : DFN1
      port map(D => N_512, CLK => HCLK_c, Q => 
        \AddressSave[4]_net_1\);
    
    \AddressSave[14]\ : DFN1
      port map(D => N_221, CLK => HCLK_c, Q => 
        \AddressSave[14]_net_1\);
    
    \Address_RNO[0]\ : OA1B
      port map(A => \haddr_c[0]\, B => N_556_i, C => 
        \Address_0_i_1[0]\, Y => N_112);
    
    ActivePhase : DFN1
      port map(D => N_108, CLK => HCLK_c, Q => \ActivePhase\);
    
    ReAddrPhase_RNO_0 : MX2
      port map(A => \ReAddrPhase\, B => N_53, S => N_48, Y => 
        N_325);
    
    \AddressSave[7]\ : DFN1
      port map(D => N_217, CLK => HCLK_c, Q => 
        \AddressSave[7]_net_1\);
    
    DataPhase_RNI0SGJ : OR3B
      port map(A => HRESETn_c, B => N_737, C => AHB_Master_In_c_3, 
        Y => N_189);
    
    \Address_RNO_0[2]\ : AO1D
      port map(A => N_949, B => N_753, C => \Address_0_i_0[2]\, Y
         => \Address_0_i_1[2]\);
    
    \AddressSave_RNO_0[22]\ : MX2
      port map(A => \AddressSave[22]_net_1\, B => N_604, S => 
        hsize_0_sqmuxa, Y => N_352);
    
    un1_AddressSave_0_sqmuxa_1_m14 : NOR3C
      port map(A => \haddr_c[12]\, B => N_13_0, C => 
        \haddr_c[13]\, Y => N_15_0);
    
    \Address_RNO[3]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[4]\, C => 
        \Address_0_i_1[3]\, Y => N_118);
    
    \Address[3]\ : DFN1
      port map(D => N_118, CLK => HCLK_c, Q => \haddr_c[3]\);
    
    \AddressSave_RNO_1[6]\ : MX2
      port map(A => N_953, B => \haddr_c[6]\, S => 
        \AddressPhase_0\, Y => N_588);
    
    ActivePhase_RNO_1 : NOR3A
      port map(A => un7_dmain(66), B => 
        ActivePhase_1_sqmuxa_i_a5_0, C => N_559, Y => N_639);
    
    un1_AddressSave_0_sqmuxa_1_m32 : XOR2
      port map(A => N_32_0, B => \haddr_c[24]\, Y => N_33_0);
    
    ReDataPhase_RNILM59 : OR2
      port map(A => \ReDataPhase\, B => \ReAddrPhase\, Y => N_559);
    
    \AddressSave_RNO_0[20]\ : MX2
      port map(A => \AddressSave[20]_net_1\, B => N_602, S => 
        hsize_0_sqmuxa, Y => N_350);
    
    \AddressSave_RNO[0]\ : NOR2B
      port map(A => N_330, B => HRESETn_c, Y => N_213);
    
    \Address_RNO_1[2]\ : OAI1
      port map(A => \AddressSave[2]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[2]\);
    
    DataPhase_RNISED9 : OR2A
      port map(A => \DataPhase\, B => AHB_Master_In_c_3, Y => 
        N_760);
    
    \Address_RNO[30]\ : OA1B
      port map(A => N_556_i, B => N_42, C => \Address_0_i_1[30]\, 
        Y => N_28);
    
    \AddressSave[0]\ : DFN1
      port map(D => N_213, CLK => HCLK_c, Q => 
        \AddressSave[0]_net_1\);
    
    AddressPhase : DFN1
      port map(D => N_191, CLK => HCLK_c, Q => \AddressPhase\);
    
    BoundaryPhase_RNO_5 : MX2A
      port map(A => \ReAddrPhase\, B => \ActivePhase\, S => 
        \AddressPhase\, Y => N_567);
    
    \AHBOut.htrans_RNO_6[0]\ : AOI1
      port map(A => N_1011, B => \AddressPhase\, C => 
        \ReAddrPhase\, Y => N_562);
    
    \AddressSave_RNO_0[5]\ : MX2
      port map(A => \AddressSave[5]_net_1\, B => N_587, S => 
        hsize_0_sqmuxa_0, Y => N_335);
    
    \AddressSave_RNO[3]\ : NOR2B
      port map(A => N_333, B => HRESETn_c, Y => 
        \AddressSave_RNO[3]_net_1\);
    
    DataPhase_RNI1I7G : OR2B
      port map(A => N_576, B => AHB_Master_In_c_3, Y => OKAY);
    
    ReAddrPhase_RNIMLKN : OR2A
      port map(A => N_1011, B => \ReAddrPhase\, Y => 
        hwrite_2_sqmuxa_1);
    
    \AddressSave_RNO[19]\ : NOR2B
      port map(A => N_349, B => HRESETn_c, Y => N_289);
    
    un1_AddressSave_0_sqmuxa_1_m42 : XNOR2
      port map(A => N_3_0, B => \haddr_c[3]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[4]\);
    
    \Address_RNO_0[6]\ : AO1D
      port map(A => N_953, B => N_753, C => \Address_0_i_0[6]\, Y
         => \Address_0_i_1[6]\);
    
    AddressPhase_RNIN7JU_0 : OR2B
      port map(A => N_756, B => N_566, Y => hsize_0_sqmuxa);
    
    un1_AddressSave_0_sqmuxa_1_m6 : OR3B
      port map(A => \haddr_c[5]\, B => \haddr_c[6]\, C => N_5_0, 
        Y => N_7_0);
    
    \AddressSave_RNO_0[17]\ : MX2
      port map(A => \AddressSave[17]_net_1\, B => N_599, S => 
        hsize_0_sqmuxa, Y => N_347);
    
    \Address[7]\ : DFN1
      port map(D => N_126, CLK => HCLK_c, Q => \haddr_c[7]\);
    
    un1_AddressSave_0_sqmuxa_1_m1 : XNOR2
      port map(A => N_566, B => \haddr_c[2]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[3]\);
    
    \Address_RNO_0[28]\ : AO1A
      port map(A => N_753_0, B => N_975, C => \Address_0_i_0[28]\, 
        Y => \Address_0_i_1[28]\);
    
    AddressPhase_RNIORDS_0 : OR2A
      port map(A => N_555, B => N_557, Y => N_753_0);
    
    \AddressSave_RNO[27]\ : NOR2B
      port map(A => N_357, B => HRESETn_c, Y => N_261);
    
    \AddressSave_RNO[12]\ : NOR2B
      port map(A => N_342, B => HRESETn_c, Y => N_285);
    
    \AddressSave[26]\ : DFN1
      port map(D => N_293, CLK => HCLK_c, Q => 
        \AddressSave[26]_net_1\);
    
    un1_AddressSave_0_sqmuxa_1_m54 : AX1C
      port map(A => \haddr_c[22]\, B => N_29_0, C => 
        \haddr_c[23]\, Y => N_55_0);
    
    un1_AddressSave_0_sqmuxa_1_m53 : XOR2
      port map(A => N_26_0, B => \haddr_c[20]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[21]\);
    
    AddressPhase_RNIORDS : OR2A
      port map(A => N_555, B => N_557, Y => N_753);
    
    \DMAOut.Ready\ : DFN1
      port map(D => N_196, CLK => HCLK_c, Q => Ready);
    
    \AddressSave[18]\ : DFN1
      port map(D => N_524, CLK => HCLK_c, Q => 
        \AddressSave[18]_net_1\);
    
    \AddressSave_RNO[30]\ : NOR2B
      port map(A => N_360, B => HRESETn_c, Y => N_532);
    
    \AddressSave_RNO[13]\ : NOR2B
      port map(A => N_343, B => HRESETn_c, Y => N_219);
    
    un1_AddressSave_0_sqmuxa_1_m29 : XOR2
      port map(A => N_29_0, B => \haddr_c[22]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[23]\);
    
    un1_AddressSave_0_sqmuxa_1_m38 : NOR3C
      port map(A => \haddr_c[26]\, B => N_36, C => \haddr_c[27]\, 
        Y => N_39);
    
    \AHBOut.hsize_RNO_0[1]\ : NOR2A
      port map(A => AHB_Master_In_c_0, B => N_554, Y => N_569);
    
    \Address_RNO_0[26]\ : AO1A
      port map(A => N_753_0, B => N_973, C => \Address_0_i_0[26]\, 
        Y => \Address_0_i_1[26]\);
    
    WriteAcc : DFN1
      port map(D => N_106, CLK => HCLK_c, Q => \WriteAcc\);
    
    \AHBOut.hsize_RNO_0[0]\ : NOR2B
      port map(A => HRESETn_c, B => \hsize_c[0]\, Y => 
        \hsize_1_i_0[0]\);
    
    EarlyPhase_RNO_0 : MX2A
      port map(A => AHB_Master_In_c_0, B => \EarlyPhase\, S => 
        un1_ahbin_3, Y => N_327);
    
    \AddressSave_RNO_0[3]\ : MX2
      port map(A => \AddressSave[3]_net_1\, B => N_595, S => 
        hsize_0_sqmuxa_0, Y => N_333);
    
    ActivePhase_RNI8O09 : OR2A
      port map(A => \ActivePhase\, B => un7_dmain(66), Y => N_560);
    
    \Address_RNO_0[29]\ : AO1D
      port map(A => N_976, B => N_753_0, C => \Address_0_i_0[29]\, 
        Y => \Address_0_i_1[29]\);
    
    un1_AddressSave_0_sqmuxa_1_m56 : XOR2
      port map(A => N_39, B => \haddr_c[28]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[29]\);
    
    un1_AddressSave_0_sqmuxa_1_m25 : NOR3C
      port map(A => \haddr_c[18]\, B => N_22_0, C => 
        \haddr_c[19]\, Y => N_26_0);
    
    un1_AddressSave_0_sqmuxa_1_m48 : XNOR2
      port map(A => N_7_0, B => \haddr_c[7]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[8]\);
    
    un1_AddressSave_0_sqmuxa_1_m20 : AX1C
      port map(A => \haddr_c[16]\, B => N_18_0, C => 
        \haddr_c[17]\, Y => \un1_AddressSave_0_sqmuxa_1_i_i[18]\);
    
    EarlyPhase_RNO_2 : OR2A
      port map(A => \ActivePhase\, B => N_761, Y => N_568);
    
    \AHBOut.htrans_RNO_1[0]\ : OR3B
      port map(A => \htrans_12_i_o2_2_4[0]\, B => 
        \htrans_12_i_o2_2_5[0]\, C => N_562, Y => 
        \htrans_RNO_1[0]\);
    
    \Address_RNO[22]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[23]\, C => 
        \Address_0_i_1[22]\, Y => N_171);
    
    \Address[9]\ : DFN1
      port map(D => N_26, CLK => HCLK_c, Q => \haddr_c[9]\);
    
    DataPhase_RNO : OA1C
      port map(A => AHB_Master_In_c_3, B => \AddressPhase_0\, C
         => DataPhase_2_i_0, Y => N_20);
    
    \Address_RNO[18]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[19]\, C => 
        \Address_0_i_1[18]\, Y => N_163);
    
    \Address_RNO_0[18]\ : AO1D
      port map(A => N_965, B => N_753_0, C => \Address_0_i_0[18]\, 
        Y => \Address_0_i_1[18]\);
    
    \AddressSave_RNO_0[28]\ : MX2
      port map(A => \AddressSave[28]_net_1\, B => N_610, S => 
        hsize_0_sqmuxa, Y => N_358);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Address_RNO[7]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[8]\, C => 
        \Address_0_i_1[7]\, Y => N_126);
    
    \Address_RNO_1[28]\ : OAI1
      port map(A => \AddressSave[28]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[28]\);
    
    \Address_RNO_0[7]\ : AO1D
      port map(A => N_954, B => N_753, C => \Address_0_i_0[7]\, Y
         => \Address_0_i_1[7]\);
    
    SingleAcc : DFN1
      port map(D => N_104, CLK => HCLK_c, Q => \SingleAcc\);
    
    \AddressSave_RNO_0[4]\ : MX2
      port map(A => \AddressSave[4]_net_1\, B => N_586, S => 
        hsize_0_sqmuxa_0, Y => N_334);
    
    \Address_RNO_1[18]\ : OAI1
      port map(A => \AddressSave[18]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[18]\);
    
    \Address[6]\ : DFN1
      port map(D => N_124, CLK => HCLK_c, Q => \haddr_c[6]\);
    
    \AddressSave_RNO_1[30]\ : MX2
      port map(A => N_977, B => \haddr_c[30]\, S => 
        \AddressPhase\, Y => N_612);
    
    \AddressSave_RNO[9]\ : NOR2B
      port map(A => N_339, B => HRESETn_c, Y => N_514);
    
    EarlyPhase_RNO_3 : AOI1B
      port map(A => N_561, B => AHB_Master_In_c_0, C => 
        AHB_Master_In_c_3, Y => un1_ahbin_3_0_0);
    
    \Address_RNO_0[16]\ : AO1D
      port map(A => N_963, B => N_753, C => \Address_0_i_0[16]\, 
        Y => \Address_0_i_1[16]\);
    
    \AddressSave_RNO_1[0]\ : MX2
      port map(A => N_947, B => \haddr_c[0]\, S => 
        \AddressPhase_0\, Y => N_592);
    
    \Address_RNO[8]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[9]\, C => 
        \Address_0_i_1[8]\, Y => N_153);
    
    \AddressSave_RNO_0[24]\ : MX2
      port map(A => \AddressSave[24]_net_1\, B => N_606, S => 
        hsize_0_sqmuxa, Y => N_354);
    
    \AddressSave[21]\ : DFN1
      port map(D => N_259, CLK => HCLK_c, Q => 
        \AddressSave[21]_net_1\);
    
    \Address_RNO_1[26]\ : OAI1
      port map(A => \AddressSave[26]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[26]\);
    
    \AddressSave_RNO_0[9]\ : MX2
      port map(A => \AddressSave[9]_net_1\, B => N_590, S => 
        hsize_0_sqmuxa_0, Y => N_339);
    
    un1_AddressSave_0_sqmuxa_1_m17 : NOR3C
      port map(A => \haddr_c[14]\, B => N_15_0, C => 
        \haddr_c[15]\, Y => N_18_0);
    
    \AHBOut.htrans_RNO_2[0]\ : AO1D
      port map(A => N_560, B => \EarlyPhase\, C => \ReAddrPhase\, 
        Y => N_676);
    
    \AddressSave_RNO_0[23]\ : MX2
      port map(A => \AddressSave[23]_net_1\, B => N_605, S => 
        hsize_0_sqmuxa, Y => N_353);
    
    SingleAcc_RNO_0 : MX2
      port map(A => \SingleAcc\, B => SingleAcc_2_sqmuxa, S => 
        hwrite_2_sqmuxa, Y => N_322);
    
    ReAddrPhase_RNI7EMV : NOR2
      port map(A => N_557, B => hwrite_2_sqmuxa_1, Y => Grant);
    
    \Address_RNO_1[16]\ : OAI1
      port map(A => \AddressSave[16]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[16]\);
    
    \Address_RNO_0[19]\ : AO1D
      port map(A => N_966, B => N_753_0, C => \Address_0_i_0[19]\, 
        Y => \Address_0_i_1[19]\);
    
    \Address[11]\ : DFN1
      port map(D => \Address_RNO[11]_net_1\, CLK => HCLK_c, Q => 
        \haddr_c[11]\);
    
    \AddressSave[31]\ : DFN1
      port map(D => N_534, CLK => HCLK_c, Q => 
        \AddressSave[31]_net_1\);
    
    \Address[31]\ : DFN1
      port map(D => N_30, CLK => HCLK_c, Q => \haddr_c[31]\);
    
    \Address_RNO_1[29]\ : OAI1
      port map(A => \AddressSave[29]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[29]\);
    
    \AddressSave_RNO_0[2]\ : MX2
      port map(A => \AddressSave[2]_net_1\, B => N_594, S => 
        hsize_0_sqmuxa_0, Y => N_332);
    
    \AddressSave[13]\ : DFN1
      port map(D => N_219, CLK => HCLK_c, Q => 
        \AddressSave[13]_net_1\);
    
    AddressPhase_RNI73CK : NOR2
      port map(A => N_554, B => \AddressPhase\, Y => N_555);
    
    DataPhase_RNI1I7G_0 : OR2A
      port map(A => Fault_0_a5_0, B => N_760, Y => Fault);
    
    \Address_RNO_1[19]\ : OAI1
      port map(A => \AddressSave[19]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[19]\);
    
    \AHBOut.hwrite_RNO_1\ : AO1B
      port map(A => N_1012, B => N_560, C => N_561, Y => N_679);
    
    \Address_RNO[2]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[3]\, C => 
        \Address_0_i_1[2]\, Y => N_116);
    
    EarlyPhase_RNI6DT61 : OA1C
      port map(A => N_561, B => N_1011, C => \un1_dmain_20_i_0\, 
        Y => N_193);
    
    \Address_RNO_1[5]\ : OAI1
      port map(A => \AddressSave[5]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[5]\);
    
    \Address_RNO[4]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[5]\, C => 
        \Address_0_i_1[4]\, Y => N_120);
    
    \AddressSave_RNO[14]\ : NOR2B
      port map(A => N_344, B => HRESETn_c, Y => N_221);
    
    EarlyPhase_RNO : NOR2B
      port map(A => N_327, B => HRESETn_c, Y => N_24);
    
    EarlyPhase_RNIHDVB : OR2
      port map(A => N_557, B => \EarlyPhase\, Y => N_758);
    
    \Address_RNO[25]\ : OA1B
      port map(A => N_556_i_0, B => N_35, C => 
        \Address_0_i_1[25]\, Y => N_177);
    
    \Address[21]\ : DFN1
      port map(D => N_169, CLK => HCLK_c, Q => \haddr_c[21]\);
    
    \AddressSave_RNO[28]\ : NOR2B
      port map(A => N_358, B => HRESETn_c, Y => N_263);
    
    \AddressSave_RNO_1[12]\ : MX2
      port map(A => N_959, B => \haddr_c[12]\, S => 
        \AddressPhase\, Y => N_617);
    
    \AddressSave_RNO_1[10]\ : MX2
      port map(A => N_957, B => \haddr_c[10]\, S => 
        \AddressPhase\, Y => N_615);
    
    ReDataPhase_RNO : NOR2B
      port map(A => N_329, B => HRESETn_c, Y => N_22);
    
    \AHBOut.hsize_RNO[0]\ : NOR2A
      port map(A => \hsize_1_i_0[0]\, B => hsize_0_sqmuxa_0, Y
         => N_149);
    
    \AddressSave_RNO[21]\ : NOR2B
      port map(A => N_351, B => HRESETn_c, Y => N_259);
    
    IdlePhase_RNO_0 : MX2B
      port map(A => \IdlePhase\, B => N_760, S => N_189, Y => 
        N_326);
    
    un1_AddressSave_0_sqmuxa_1_m57 : AX1C
      port map(A => \haddr_c[28]\, B => N_39, C => \haddr_c[29]\, 
        Y => N_58_0);
    
    \Address[17]\ : DFN1
      port map(D => N_161, CLK => HCLK_c, Q => \haddr_c[17]\);
    
    \AddressSave[10]\ : DFN1
      port map(D => N_516, CLK => HCLK_c, Q => 
        \AddressSave[10]_net_1\);
    
    \AddressSave_RNO_0[26]\ : MX2
      port map(A => \AddressSave[26]_net_1\, B => N_608, S => 
        hsize_0_sqmuxa, Y => N_356);
    
    \Address_RNO_1[1]\ : OAI1
      port map(A => \AddressSave[1]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[1]\);
    
    \Address_RNO_1[6]\ : OAI1
      port map(A => \AddressSave[6]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[6]\);
    
    un1_AddressSave_0_sqmuxa_1_m51 : AX1C
      port map(A => \haddr_c[12]\, B => N_13_0, C => 
        \haddr_c[13]\, Y => \un1_AddressSave_0_sqmuxa_1_i_i[14]\);
    
    un1_AddressSave_0_sqmuxa_1_m34 : AX1C
      port map(A => \haddr_c[24]\, B => N_32_0, C => 
        \haddr_c[25]\, Y => N_35);
    
    \Address_RNIV6FD[9]\ : NOR2B
      port map(A => \haddr_c[9]\, B => \haddr_c[2]\, Y => 
        \htrans_12_i_o2_2_0[0]\);
    
    \Address[27]\ : DFN1
      port map(D => N_128, CLK => HCLK_c, Q => \haddr_c[27]\);
    
    \AddressSave[3]\ : DFN1
      port map(D => \AddressSave_RNO[3]_net_1\, CLK => HCLK_c, Q
         => \AddressSave[3]_net_1\);
    
    DataPhase : DFN1
      port map(D => N_20, CLK => HCLK_c, Q => \DataPhase\);
    
    \AddressSave[2]\ : DFN1
      port map(D => \AddressSave_RNO[2]_net_1\, CLK => HCLK_c, Q
         => \AddressSave[2]_net_1\);
    
    \AddressSave[27]\ : DFN1
      port map(D => N_261, CLK => HCLK_c, Q => 
        \AddressSave[27]_net_1\);
    
    AddressPhase_0 : DFN1
      port map(D => N_191, CLK => HCLK_c, Q => \AddressPhase_0\);
    
    \Address_RNO_0[20]\ : AO1D
      port map(A => N_967, B => N_753_0, C => \Address_0_i_0[20]\, 
        Y => \Address_0_i_1[20]\);
    
    \AddressSave_RNO[8]\ : NOR2B
      port map(A => N_338, B => HRESETn_c, Y => N_283);
    
    \AddressSave[5]\ : DFN1
      port map(D => N_281, CLK => HCLK_c, Q => 
        \AddressSave[5]_net_1\);
    
    \AddressSave[24]\ : DFN1
      port map(D => N_528, CLK => HCLK_c, Q => 
        \AddressSave[24]_net_1\);
    
    \AddressSave_RNO_1[8]\ : MX2
      port map(A => N_955, B => \haddr_c[8]\, S => \AddressPhase\, 
        Y => N_613);
    
    \Address_RNO[31]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[32]\, C => 
        \Address_0_i_1[31]\, Y => N_30);
    
    \AHBOut.htrans_RNO_4[0]\ : OR2A
      port map(A => \ReAddrPhase\, B => \AddressPhase\, Y => 
        N_678);
    
    \AHBOut.htrans_RNO[0]\ : NOR3C
      port map(A => \htrans_12_i_2[0]\, B => \htrans_RNO_1[0]\, C
         => N_676, Y => N_137_i_0);
    
    un1_AddressSave_0_sqmuxa_1_m44 : XNOR2
      port map(A => N_5_0, B => \haddr_c[5]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[6]\);
    
    un1_AddressSave_0_sqmuxa_1_m43 : AX1
      port map(A => N_3_0, B => \haddr_c[3]\, C => \haddr_c[4]\, 
        Y => \un1_AddressSave_0_sqmuxa_1_i_i[5]\);
    
    \Address_RNO[12]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[13]\, C => 
        \Address_0_i_1[12]\, Y => \Address_RNO[12]_net_1\);
    
    DataPhase_RNIGGQC_0 : NOR2A
      port map(A => \DataPhase\, B => N_558, Y => N_576);
    
    un1_AddressSave_0_sqmuxa_1_m36 : XOR2
      port map(A => N_36, B => \haddr_c[26]\, Y => N_37);
    
    \Address_RNO_0[23]\ : AO1D
      port map(A => N_970, B => N_753_0, C => \Address_0_i_0[23]\, 
        Y => \Address_0_i_1[23]\);
    
    un1_AddressSave_0_sqmuxa_1_m22 : XOR2
      port map(A => N_22_0, B => \haddr_c[18]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[19]\);
    
    \AddressSave_RNO[6]\ : NOR2B
      port map(A => N_336, B => HRESETn_c, Y => N_215);
    
    \AddressSave_RNO_0[29]\ : MX2
      port map(A => \AddressSave[29]_net_1\, B => N_611, S => 
        hsize_0_sqmuxa, Y => N_359);
    
    \Address[1]\ : DFN1
      port map(D => N_114, CLK => HCLK_c, Q => \haddr_c[1]\);
    
    \AddressSave_RNO[20]\ : NOR2B
      port map(A => N_350, B => HRESETn_c, Y => N_225);
    
    \AddressSave_RNO[17]\ : NOR2B
      port map(A => N_347, B => HRESETn_c, Y => N_522);
    
    un1_AddressSave_0_sqmuxa_1_m46 : AX1
      port map(A => N_7_0, B => \haddr_c[7]\, C => \haddr_c[8]\, 
        Y => \un1_AddressSave_0_sqmuxa_1_i_i[9]\);
    
    \AHBOut.hburst[1]\ : DFN1E1
      port map(D => N_682, CLK => HCLK_c, E => N_130, Q => 
        hburst_c(1));
    
    ReDataPhase_RNIHO18_0 : OR2A
      port map(A => \ReDataPhase\, B => N_553, Y => N_754_0);
    
    un1_dmain_20_i_0 : OR2A
      port map(A => HRESETn_c, B => N_553, Y => 
        \un1_dmain_20_i_0\);
    
    un1_AddressSave_0_sqmuxa_1_m4 : OR3B
      port map(A => \haddr_c[3]\, B => \haddr_c[4]\, C => N_3_0, 
        Y => N_5_0);
    
    ReAddrPhase_RNI25HF : NOR3A
      port map(A => HRESETn_c, B => \ReAddrPhase\, C => 
        time_select_0, Y => \hburst_11_i_a2_i_a5_1[1]\);
    
    AddressPhase_RNIN7JU : OR2B
      port map(A => N_756, B => N_566, Y => hsize_0_sqmuxa_0);
    
    BoundaryPhase_RNO_4 : OR3C
      port map(A => N_829, B => N_567, C => N_1011, Y => N_684);
    
    \AddressSave_RNO_1[18]\ : MX2
      port map(A => N_965, B => \haddr_c[18]\, S => 
        \AddressPhase_0\, Y => N_600);
    
    \AddressSave_RNO_0[25]\ : MX2
      port map(A => \AddressSave[25]_net_1\, B => N_607, S => 
        hsize_0_sqmuxa, Y => N_355);
    
    AddressPhase_RNIKTLA : MX2C
      port map(A => \AddressPhase\, B => AHB_Master_In_c_0, S => 
        AHB_Master_In_c_3, Y => N_614);
    
    \AddressSave_RNO_0[21]\ : MX2
      port map(A => \AddressSave[21]_net_1\, B => N_603, S => 
        hsize_0_sqmuxa, Y => N_351);
    
    \Address_RNO_0[10]\ : AO1D
      port map(A => N_957, B => N_753, C => \Address_0_i_0[10]\, 
        Y => \Address_0_i_1[10]\);
    
    \Address_RNO[20]\ : OA1B
      port map(A => N_556_i_0, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[21]\, C => 
        \Address_0_i_1[20]\, Y => N_167);
    
    ActivePhase_RNO_0 : AO1A
      port map(A => N_639, B => \ActivePhase\, C => 
        hwrite_2_sqmuxa, Y => N_320);
    
    \AddressSave_RNO[26]\ : NOR2B
      port map(A => N_356, B => HRESETn_c, Y => N_293);
    
    \Address_RNO_1[20]\ : OAI1
      port map(A => \AddressSave[20]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[20]\);
    
    \AHBOut.htrans_RNO_3[0]\ : NOR2A
      port map(A => HRESETn_c, B => N_557, Y => 
        \htrans_12_i_0[0]\);
    
    \AddressSave[28]\ : DFN1
      port map(D => N_263, CLK => HCLK_c, Q => 
        \AddressSave[28]_net_1\);
    
    ReDataPhase_RNIHO18_1 : OR2
      port map(A => \ReDataPhase\, B => N_553, Y => N_557);
    
    \AddressSave_RNO_1[4]\ : MX2
      port map(A => N_951, B => \haddr_c[4]\, S => 
        \AddressPhase_0\, Y => N_586);
    
    EarlyPhase_RNIFRKC1 : NOR3A
      port map(A => N_560, B => hwrite_2_sqmuxa_1, C => N_758, Y
         => hwrite_2_sqmuxa);
    
    \Address_RNO_1[10]\ : OAI1
      port map(A => \AddressSave[10]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[10]\);
    
    \AddressSave_RNO_1[22]\ : MX2
      port map(A => N_969, B => \haddr_c[22]\, S => 
        \AddressPhase_0\, Y => N_604);
    
    \Address_RNI2O5T1[4]\ : NOR3B
      port map(A => \htrans_12_i_o2_2_4[0]\, B => 
        \htrans_12_i_o2_2_5[0]\, C => N_566, Y => N_580);
    
    ReDataPhase : DFN1
      port map(D => N_22, CLK => HCLK_c, Q => \ReDataPhase\);
    
    \AHBOut.htrans[0]\ : DFN1E1
      port map(D => N_137_i_0, CLK => HCLK_c, E => N_189, Q => 
        htrans_c(0));
    
    EarlyPhase_RNIQH6K : NOR2
      port map(A => un7_dmain(66), B => N_758, Y => N_829);
    
    BoundaryPhase_RNO_3 : OR3B
      port map(A => \ReAddrPhase\, B => \AddressPhase\, C => 
        N_557, Y => N_686);
    
    un1_AddressSave_0_sqmuxa_1_m15 : XOR2
      port map(A => N_15_0, B => \haddr_c[14]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[15]\);
    
    ReDataPhase_RNO_0 : AO1
      port map(A => \ReDataPhase\, B => N_553, C => Retry, Y => 
        N_329);
    
    \AddressSave_RNO_1[20]\ : MX2
      port map(A => N_967, B => \haddr_c[20]\, S => 
        \AddressPhase_0\, Y => N_602);
    
    \AddressSave_RNO_1[14]\ : MX2
      port map(A => N_961, B => \haddr_c[14]\, S => 
        \AddressPhase_0\, Y => N_596);
    
    un1_AddressSave_0_sqmuxa_1_m8 : OR3B
      port map(A => \haddr_c[7]\, B => \haddr_c[8]\, C => N_7_0, 
        Y => N_9_0);
    
    un1_AddressSave_0_sqmuxa_1_m28 : NOR3C
      port map(A => \haddr_c[20]\, B => N_26_0, C => 
        \haddr_c[21]\, Y => N_29_0);
    
    \Address_RNO_0[13]\ : AO1D
      port map(A => N_960, B => N_753, C => \Address_0_i_0[13]\, 
        Y => \Address_0_i_1[13]\);
    
    \Address_RNO[15]\ : OA1B
      port map(A => N_556_i, B => 
        \un1_AddressSave_0_sqmuxa_1_i_i[16]\, C => 
        \Address_0_i_1[15]\, Y => N_157);
    
    ActivePhase_RNIB5HP : OR3B
      port map(A => AHB_Master_In_c_0, B => N_561, C => N_560, Y
         => N_582);
    
    un1_AddressSave_0_sqmuxa_1_m10 : XOR2
      port map(A => N_580, B => \haddr_c[10]\, Y => 
        \un1_AddressSave_0_sqmuxa_1_i_i[11]\);
    
    \AHBOut.hburst_RNO[0]\ : OA1A
      port map(A => N_561, B => N_1011, C => 
        \hburst_11_0_a2_i_2[0]\, Y => N_56_i_0);
    
    \AddressSave_RNO_1[13]\ : MX2
      port map(A => N_960, B => \haddr_c[13]\, S => 
        \AddressPhase\, Y => N_618);
    
    \Address_RNO_1[23]\ : OAI1
      port map(A => \AddressSave[23]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[23]\);
    
    \Address_RNO_0[21]\ : AO1D
      port map(A => N_968, B => N_753_0, C => \Address_0_i_0[21]\, 
        Y => \Address_0_i_1[21]\);
    
    \AddressSave[19]\ : DFN1
      port map(D => N_289, CLK => HCLK_c, Q => 
        \AddressSave[19]_net_1\);
    
    ReDataPhase_RNI5AUG : NOR2
      port map(A => N_1011, B => \ReDataPhase\, Y => N_635);
    
    \Address_RNO_1[13]\ : OAI1
      port map(A => \AddressSave[13]_net_1\, B => N_754, C => 
        HRESETn_c, Y => \Address_0_i_0[13]\);
    
    un1_AddressSave_0_sqmuxa_1_m59 : AX1C
      port map(A => \haddr_c[30]\, B => N_41, C => \haddr_c[31]\, 
        Y => \un1_AddressSave_0_sqmuxa_1_i_i[32]\);
    
    \Address_RNO_1[9]\ : OAI1
      port map(A => \AddressSave[9]_net_1\, B => N_754_0, C => 
        HRESETn_c, Y => \Address_0_i_0[9]\);
    
    \Address_RNO_0[0]\ : AO1D
      port map(A => N_947, B => N_753_0, C => \Address_0_i_0[0]\, 
        Y => \Address_0_i_1[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_dma is

    port( addr_data_f0       : in    std_logic_vector(31 downto 0);
          addr_data_f1       : in    std_logic_vector(31 downto 0);
          addr_data_f2       : in    std_logic_vector(31 downto 0);
          addr_data_f3       : in    std_logic_vector(31 downto 0);
          status_full        : out   std_logic_vector(3 downto 0);
          status_full_err    : out   std_logic_vector(3 downto 0);
          nb_burst_available : in    std_logic_vector(10 downto 0);
          haddr_c            : out   std_logic_vector(31 downto 0);
          AHB_Master_In_c_3  : in    std_logic;
          AHB_Master_In_c_0  : in    std_logic;
          AHB_Master_In_c_4  : in    std_logic;
          AHB_Master_In_c_5  : in    std_logic;
          hsize_c            : out   std_logic_vector(1 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          hburst_c           : out   std_logic_vector(2 downto 0);
          status_full_ack    : in    std_logic_vector(3 downto 0);
          ready_i_0          : in    std_logic_vector(3 downto 0);
          data_ren           : out   std_logic_vector(3 downto 0);
          time_ren           : out   std_logic_vector(3 downto 0);
          time_ren_1z        : out   std_logic;
          data_ren_1z        : out   std_logic;
          N_43               : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          hwrite_c           : out   std_logic;
          un20_time_write    : out   std_logic;
          un13_time_write    : out   std_logic;
          HRESETn_c          : in    std_logic;
          HCLK_c             : in    std_logic
        );

end lpp_waveform_dma;

architecture DEF_ARCH of lpp_waveform_dma is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\
    port( nb_burst_available  : in    std_logic_vector(10 downto 0) := (others => 'U');
          status_full_err     : out   std_logic_vector(2 to 2);
          status_full         : out   std_logic_vector(2 to 2);
          sel_data            : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_1          : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_0          : in    std_logic_vector(1 to 1) := (others => 'U');
          update_and_sel_3    : in    std_logic_vector(5 downto 4) := (others => 'U');
          addr_data_f2        : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full_ack     : in    std_logic_vector(2 to 2) := (others => 'U');
          addr_data_vector_62 : out   std_logic;
          addr_data_vector_61 : out   std_logic;
          addr_data_vector_5  : in    std_logic := 'U';
          addr_data_vector_4  : in    std_logic := 'U';
          addr_data_vector_3  : in    std_logic := 'U';
          addr_data_vector_0  : in    std_logic := 'U';
          addr_data_vector_12 : in    std_logic := 'U';
          addr_data_vector_11 : in    std_logic := 'U';
          addr_data_vector_9  : in    std_logic := 'U';
          addr_data_vector_7  : in    std_logic := 'U';
          addr_data_vector_6  : in    std_logic := 'U';
          addr_data_vector_26 : in    std_logic := 'U';
          addr_data_vector_24 : in    std_logic := 'U';
          addr_data_vector_22 : in    std_logic := 'U';
          addr_data_vector_28 : in    std_logic := 'U';
          addr_data_vector_66 : out   std_logic;
          addr_data_vector_65 : out   std_logic;
          addr_data_vector_91 : out   std_logic;
          addr_data_vector_89 : out   std_logic;
          addr_data_vector_87 : out   std_logic;
          addr_data_vector_63 : out   std_logic;
          addr_data_vector_72 : out   std_logic;
          addr_data_vector_74 : out   std_logic;
          addr_data_vector_79 : out   std_logic;
          addr_data_vector_78 : out   std_logic;
          addr_data_vector_81 : out   std_logic;
          addr_data_vector_80 : out   std_logic;
          addr_data_vector_84 : out   std_logic;
          addr_data_vector_85 : out   std_logic;
          addr_data_vector_77 : out   std_logic;
          addr_data_vector_82 : out   std_logic;
          addr_data_vector_83 : out   std_logic;
          N_1329              : out   std_logic;
          N_1328              : out   std_logic;
          N_1327              : out   std_logic;
          N_1324              : out   std_logic;
          N_1322              : out   std_logic;
          N_1321              : out   std_logic;
          N_1319              : out   std_logic;
          N_1317              : out   std_logic;
          N_1316              : out   std_logic;
          N_1308              : out   std_logic;
          N_1306              : out   std_logic;
          N_1304              : out   std_logic;
          N_1296              : out   std_logic;
          HRESETn_c           : in    std_logic := 'U';
          HCLK_c              : in    std_logic := 'U'
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\
    port( nb_burst_available  : in    std_logic_vector(10 downto 0) := (others => 'U');
          status_full_err     : out   std_logic_vector(0 to 0);
          status_full         : out   std_logic_vector(0 to 0);
          sel_data            : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_1          : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_0          : in    std_logic_vector(1 to 1) := (others => 'U');
          update_and_sel_7    : in    std_logic_vector(1 downto 0) := (others => 'U');
          addr_data_f0        : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full_ack     : in    std_logic_vector(0 to 0) := (others => 'U');
          addr_data_vector_69 : in    std_logic := 'U';
          addr_data_vector_68 : in    std_logic := 'U';
          addr_data_vector_66 : in    std_logic := 'U';
          addr_data_vector_77 : in    std_logic := 'U';
          addr_data_vector_75 : in    std_logic := 'U';
          addr_data_vector_86 : in    std_logic := 'U';
          addr_data_vector_85 : in    std_logic := 'U';
          addr_data_vector_84 : in    std_logic := 'U';
          addr_data_vector_83 : in    std_logic := 'U';
          addr_data_vector_82 : in    std_logic := 'U';
          addr_data_vector_81 : in    std_logic := 'U';
          addr_data_vector_80 : in    std_logic := 'U';
          addr_data_vector_92 : in    std_logic := 'U';
          addr_data_vector_90 : in    std_logic := 'U';
          addr_data_vector_88 : in    std_logic := 'U';
          addr_data_vector_87 : in    std_logic := 'U';
          addr_data_vector_94 : in    std_logic := 'U';
          addr_data_vector_65 : in    std_logic := 'U';
          addr_data_vector_64 : in    std_logic := 'U';
          addr_data_vector_3  : out   std_logic;
          addr_data_vector_31 : out   std_logic;
          addr_data_vector_14 : out   std_logic;
          addr_data_vector_15 : out   std_logic;
          addr_data_vector_27 : out   std_logic;
          addr_data_vector_29 : out   std_logic;
          addr_data_vector_25 : out   std_logic;
          addr_data_vector_6  : out   std_logic;
          addr_data_vector_8  : out   std_logic;
          addr_data_vector_7  : out   std_logic;
          addr_data_vector_10 : out   std_logic;
          addr_data_vector_9  : out   std_logic;
          addr_data_vector_12 : out   std_logic;
          N_1326              : out   std_logic;
          N_1325              : out   std_logic;
          N_1323              : out   std_logic;
          N_1320              : out   std_logic;
          N_1318              : out   std_logic;
          N_1315              : out   std_logic;
          N_1314              : out   std_logic;
          N_1313              : out   std_logic;
          N_1312              : out   std_logic;
          N_1311              : out   std_logic;
          N_1310              : out   std_logic;
          N_1309              : out   std_logic;
          N_1307              : out   std_logic;
          N_1305              : out   std_logic;
          N_1303              : out   std_logic;
          N_1302              : out   std_logic;
          N_1295              : out   std_logic;
          N_1280              : out   std_logic;
          N_1279              : out   std_logic;
          HRESETn_c           : in    std_logic := 'U';
          HCLK_c              : in    std_logic := 'U'
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component lpp_dma_send_16word
    port( un7_dmain        : out   std_logic_vector(66 to 66);
          data_address     : in    std_logic_vector(31 downto 0) := (others => 'U');
          Store            : out   std_logic;
          Fault            : in    std_logic := 'U';
          un1_data_send_ok : out   std_logic;
          Request_0        : in    std_logic := 'U';
          N_1011           : out   std_logic;
          Lock_0           : in    std_logic := 'U';
          N_1013           : out   std_logic;
          N_957            : out   std_logic;
          N_956            : out   std_logic;
          N_955            : out   std_logic;
          N_954            : out   std_logic;
          N_953            : out   std_logic;
          N_952            : out   std_logic;
          N_951            : out   std_logic;
          N_964            : out   std_logic;
          N_963            : out   std_logic;
          N_962            : out   std_logic;
          N_961            : out   std_logic;
          N_960            : out   std_logic;
          time_select      : in    std_logic := 'U';
          N_959            : out   std_logic;
          N_958            : out   std_logic;
          N_971            : out   std_logic;
          N_970            : out   std_logic;
          N_969            : out   std_logic;
          N_968            : out   std_logic;
          N_967            : out   std_logic;
          N_966            : out   std_logic;
          N_965            : out   std_logic;
          N_978            : out   std_logic;
          N_977            : out   std_logic;
          N_976            : out   std_logic;
          N_975            : out   std_logic;
          N_974            : out   std_logic;
          N_973            : out   std_logic;
          N_972            : out   std_logic;
          N_950            : out   std_logic;
          N_949            : out   std_logic;
          N_948            : out   std_logic;
          time_select_0    : in    std_logic := 'U';
          N_947            : out   std_logic;
          N_249            : out   std_logic;
          Grant            : in    std_logic := 'U';
          Ready            : in    std_logic := 'U';
          data_send        : in    std_logic := 'U';
          OKAY             : in    std_logic := 'U';
          N_200            : out   std_logic;
          HRESETn_c        : in    std_logic := 'U';
          HCLK_c           : in    std_logic := 'U'
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\
    port( nb_burst_available  : in    std_logic_vector(10 downto 0) := (others => 'U');
          status_full_err     : out   std_logic_vector(1 to 1);
          status_full         : out   std_logic_vector(1 to 1);
          sel_data            : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_0          : in    std_logic_vector(1 to 1) := (others => 'U');
          update_and_sel_5    : in    std_logic_vector(3 downto 2) := (others => 'U');
          addr_data_f1        : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full_ack     : in    std_logic_vector(1 to 1) := (others => 'U');
          addr_data_vector_94 : in    std_logic := 'U';
          addr_data_vector_91 : in    std_logic := 'U';
          addr_data_vector_89 : in    std_logic := 'U';
          addr_data_vector_87 : in    std_logic := 'U';
          addr_data_vector_86 : in    std_logic := 'U';
          addr_data_vector_85 : in    std_logic := 'U';
          addr_data_vector_84 : in    std_logic := 'U';
          addr_data_vector_83 : in    std_logic := 'U';
          addr_data_vector_67 : in    std_logic := 'U';
          addr_data_vector_66 : in    std_logic := 'U';
          addr_data_vector_65 : in    std_logic := 'U';
          addr_data_vector_64 : in    std_logic := 'U';
          addr_data_vector_75 : in    std_logic := 'U';
          addr_data_vector_73 : in    std_logic := 'U';
          addr_data_vector_81 : in    std_logic := 'U';
          addr_data_vector_79 : in    std_logic := 'U';
          addr_data_vector_77 : in    std_logic := 'U';
          addr_data_vector_24 : out   std_logic;
          addr_data_vector_31 : out   std_logic;
          addr_data_vector_16 : out   std_logic;
          addr_data_vector_14 : out   std_logic;
          addr_data_vector_18 : out   std_logic;
          addr_data_vector_26 : out   std_logic;
          addr_data_vector_29 : out   std_logic;
          addr_data_vector_28 : out   std_logic;
          addr_data_vector_5  : out   std_logic;
          addr_data_vector_4  : out   std_logic;
          addr_data_vector_6  : out   std_logic;
          addr_data_vector_12 : out   std_logic;
          addr_data_vector_10 : out   std_logic;
          addr_data_vector_7  : out   std_logic;
          addr_data_vector_8  : out   std_logic;
          N_913               : out   std_logic;
          N_910               : out   std_logic;
          N_908               : out   std_logic;
          N_906               : out   std_logic;
          N_905               : out   std_logic;
          N_904               : out   std_logic;
          N_903               : out   std_logic;
          N_902               : out   std_logic;
          N_1300              : out   std_logic;
          N_1299              : out   std_logic;
          N_1298              : out   std_logic;
          N_1297              : out   std_logic;
          N_1294              : out   std_logic;
          N_1292              : out   std_logic;
          N_1286              : out   std_logic;
          N_1284              : out   std_logic;
          N_1282              : out   std_logic;
          HRESETn_c           : in    std_logic := 'U';
          HCLK_c              : in    std_logic := 'U'
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component lpp_dma_send_1word
    port( Lock             : out   std_logic;
          Request          : out   std_logic;
          HRESETn_c        : in    std_logic := 'U';
          HCLK_c           : in    std_logic := 'U';
          un1_time_send_ok : out   std_logic;
          time_select      : in    std_logic := 'U';
          Store            : in    std_logic := 'U';
          N_1012           : out   std_logic;
          Ready            : in    std_logic := 'U';
          Fault            : in    std_logic := 'U';
          time_send        : in    std_logic := 'U';
          Grant            : in    std_logic := 'U'
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\
    port( nb_burst_available  : in    std_logic_vector(10 downto 0) := (others => 'U');
          status_full_err     : out   std_logic_vector(3 to 3);
          status_full         : out   std_logic_vector(3 to 3);
          sel_data            : in    std_logic_vector(1 to 1) := (others => 'U');
          sel_data_0          : in    std_logic_vector(1 to 1) := (others => 'U');
          update_and_sel_1    : in    std_logic_vector(7 downto 6) := (others => 'U');
          addr_data_f3        : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full_ack     : in    std_logic_vector(3 to 3) := (others => 'U');
          addr_data_vector_61 : out   std_logic;
          addr_data_vector_60 : out   std_logic;
          addr_data_vector_27 : in    std_logic := 'U';
          addr_data_vector_25 : in    std_logic := 'U';
          addr_data_vector_24 : in    std_logic := 'U';
          addr_data_vector_22 : in    std_logic := 'U';
          addr_data_vector_20 : in    std_logic := 'U';
          addr_data_vector_0  : in    std_logic := 'U';
          addr_data_vector_6  : in    std_logic := 'U';
          addr_data_vector_4  : in    std_logic := 'U';
          addr_data_vector_3  : in    std_logic := 'U';
          addr_data_vector_2  : in    std_logic := 'U';
          addr_data_vector_1  : in    std_logic := 'U';
          addr_data_vector_14 : in    std_logic := 'U';
          addr_data_vector_12 : in    std_logic := 'U';
          addr_data_vector_10 : in    std_logic := 'U';
          addr_data_vector_8  : in    std_logic := 'U';
          addr_data_vector_63 : out   std_logic;
          addr_data_vector_90 : out   std_logic;
          addr_data_vector_87 : out   std_logic;
          addr_data_vector_85 : out   std_logic;
          addr_data_vector_62 : out   std_logic;
          addr_data_vector_69 : out   std_logic;
          addr_data_vector_73 : out   std_logic;
          addr_data_vector_71 : out   std_logic;
          addr_data_vector_77 : out   std_logic;
          addr_data_vector_79 : out   std_logic;
          addr_data_vector_82 : out   std_logic;
          addr_data_vector_83 : out   std_logic;
          addr_data_vector_75 : out   std_logic;
          addr_data_vector_80 : out   std_logic;
          addr_data_vector_81 : out   std_logic;
          N_914               : out   std_logic;
          N_912               : out   std_logic;
          N_911               : out   std_logic;
          N_909               : out   std_logic;
          N_907               : out   std_logic;
          N_1301              : out   std_logic;
          N_1293              : out   std_logic;
          N_1291              : out   std_logic;
          N_1290              : out   std_logic;
          N_1289              : out   std_logic;
          N_1288              : out   std_logic;
          N_1287              : out   std_logic;
          N_1285              : out   std_logic;
          N_1283              : out   std_logic;
          N_1281              : out   std_logic;
          HRESETn_c           : in    std_logic := 'U';
          HCLK_c              : in    std_logic := 'U'
        );
  end component;

  component DMA2AHB
    port( hburst_c           : out   std_logic_vector(2 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          un7_dmain          : in    std_logic_vector(66 to 66) := (others => 'U');
          hsize_c            : out   std_logic_vector(1 downto 0);
          AHB_Master_In_c_5  : in    std_logic := 'U';
          AHB_Master_In_c_4  : in    std_logic := 'U';
          AHB_Master_In_c_0  : in    std_logic := 'U';
          AHB_Master_In_c_3  : in    std_logic := 'U';
          haddr_c            : out   std_logic_vector(31 downto 0);
          hwrite_c           : out   std_logic;
          Ready              : out   std_logic;
          N_1012             : in    std_logic := 'U';
          Grant              : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          OKAY               : out   std_logic;
          Fault              : out   std_logic;
          N_1011             : in    std_logic := 'U';
          N_1013             : in    std_logic := 'U';
          N_43               : out   std_logic;
          time_select_0      : in    std_logic := 'U';
          N_960              : in    std_logic := 'U';
          N_959              : in    std_logic := 'U';
          N_958              : in    std_logic := 'U';
          N_957              : in    std_logic := 'U';
          N_964              : in    std_logic := 'U';
          N_963              : in    std_logic := 'U';
          N_962              : in    std_logic := 'U';
          N_961              : in    std_logic := 'U';
          N_955              : in    std_logic := 'U';
          N_954              : in    std_logic := 'U';
          N_953              : in    std_logic := 'U';
          N_952              : in    std_logic := 'U';
          N_951              : in    std_logic := 'U';
          N_950              : in    std_logic := 'U';
          N_949              : in    std_logic := 'U';
          N_948              : in    std_logic := 'U';
          N_947              : in    std_logic := 'U';
          N_956              : in    std_logic := 'U';
          N_965              : in    std_logic := 'U';
          N_966              : in    std_logic := 'U';
          N_967              : in    std_logic := 'U';
          N_968              : in    std_logic := 'U';
          N_969              : in    std_logic := 'U';
          N_970              : in    std_logic := 'U';
          N_971              : in    std_logic := 'U';
          N_972              : in    std_logic := 'U';
          N_973              : in    std_logic := 'U';
          N_974              : in    std_logic := 'U';
          N_975              : in    std_logic := 'U';
          N_976              : in    std_logic := 'U';
          N_977              : in    std_logic := 'U';
          HRESETn_c          : in    std_logic := 'U';
          N_978              : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U'
        );
  end component;

    signal count_send_time_e18_0_0, \count_send_time[18]_net_1\, 
        N_1220, N_1099, \count_send_time_RNO[17]_net_1\, N_1091, 
        N_1096, N_1137, \count_send_time_RNO[28]_net_1\, N_1156, 
        \count_send_time[28]_net_1\, 
        \count_send_time_RNO[29]_net_1\, N_1160, 
        \count_send_time[29]_net_1\, count_send_time_e31, N_1191, 
        N_1193, N_1194, count_send_time_e30, N_1126, 
        count_send_time_e30_0_0, N_1128, N_1146, 
        \count_send_time[27]_net_1\, count_send_time_e30_0_a2_2_1, 
        count_send_time_e25, N_1178, N_1177, N_1180, 
        count_send_time_e24, N_1173, N_1172, N_1175, N_1161, 
        \count_send_time[31]_net_1\, \state[2]_net_1\, N_1162, 
        N_1145_0, \count_send_time[25]_net_1\, 
        count_send_time_e25_0_o3_N_7_i_0, 
        \count_send_time[23]_net_1\, N_1069, 
        count_send_time_e24_0_a2_1_0, 
        count_send_time_e24_0_a2_0_0, count_send_time_e23, N_1121, 
        N_1122, N_1123, count_send_time_e22, N_1117, N_1118, 
        N_1119, count_send_time_e21, N_1112, N_1113, N_1114, 
        count_send_time_e20, N_1107, N_1108, N_1109, 
        count_send_time_e19, N_1103, N_1102, N_1104, 
        count_send_time_e18, count_send_time_e30_0_a2_0_0, 
        \count_send_time[21]_net_1\, N_1066, 
        count_send_time_e22_0_a2_1_0, count_send_time_e22_0_a2_0, 
        N_1145, N_1063, \count_send_time[19]_net_1\, 
        count_send_time_e20_0_a2_1_0, count_send_time_e20_0_a2_0, 
        \count_send_time[17]_net_1\, N_1061, 
        count_send_time_e18_0_a2_0_0, N_1059, 
        \count_send_time[15]_net_1\, 
        count_send_time_e25_0_o3_m6_0_a2_7, N_1057, 
        \count_send_time[11]_net_1\, \count_send_time[12]_net_1\, 
        N_1159, \count_send_time[13]_net_1\, 
        \count_send_time[14]_net_1\, \count_send_time[16]_net_1\, 
        \count_send_time[20]_net_1\, \count_send_time[22]_net_1\, 
        \count_send_time_RNO[26]_net_1\, N_1163, 
        \count_send_time[26]_net_1\, 
        \count_send_time_RNO[27]_net_1\, N_1164, 
        \count_send_time[9]_net_1\, \count_send_time[10]_net_1\, 
        N_1225, N_1217, \count_send_time[0]_net_1\, 
        \count_send_time[1]_net_1\, \count_send_time[2]_net_1\, 
        N_1219, \count_send_time[3]_net_1\, 
        \count_send_time[4]_net_1\, N_1223, 
        \count_send_time[5]_net_1\, \count_send_time[6]_net_1\, 
        \count_send_time[7]_net_1\, \count_send_time[8]_net_1\, 
        \sel_data_0[0]_net_1\, N_1016_i_0, \state[7]_net_1\, 
        \sel_data_1[1]_net_1\, N_1015, \sel_data_0[1]_net_1\, 
        \state_0[2]_net_1\, \state_ns_i_a2_0[5]_net_1\, 
        \time_select_0\, time_fifo_ren_1, N_816, 
        time_fifo_ren_1_i, N_1049, N_1026, \state[4]_net_1\, 
        \state_ns_i_a2_0_1[5]\, N_1048, \state_ns_i_a2_0_0[5]\, 
        \count_send_time[24]_net_1\, \count_send_time[30]_net_1\, 
        N_1125, N_1075, count_send_time_e16_i_0, N_1077, 
        \state_ns_i_a2_0_a4_0_19_i[5]\, N_1050, 
        count_send_time_e25_0_o3_m6_0_a2_2, 
        count_send_time_e25_0_o3_m6_0_a2_1, 
        count_send_time_e25_0_o3_m6_0_a2_6, 
        count_send_time_e25_0_o3_m6_0_a2_4, 
        count_send_time_e14_i_0, 
        \count_send_time_RNO_1[14]_net_1\, state_tr2_i_0, 
        \send_16_3_time[0]_net_1\, 
        \state_ns_i_a2_0_a3_0[5]_net_1\, 
        \send_16_3_time_1_sqmuxa_i_o3_0\, 
        count_send_time_e12_0_a2_0_0, 
        count_send_time_e12_0_a2_1_0, count_send_time_e10_0_a2_0, 
        count_send_time_e10_0_a2_1_0, count_send_time_e8_0_a2_0, 
        count_send_time_e8_0_a2_1_0, count_send_time_e2_0_a2_1_0, 
        state_tr13_0_a2_15, state_tr13_0_a2_9_0, 
        state_tr13_0_a2_8, state_tr13_0_a2_12, state_tr13_0_a2_14, 
        state_tr13_0_a2_10, state_tr13_0_a2_9, state_tr13_0_a2_7, 
        state_tr13_0_a2_17_0, state_tr13_0_a2_17_1, 
        state_tr13_0_a2_6, state_tr13_0_a2_4, state_tr13_0_a2_2, 
        \state_ns_i_a2_0_a4_0_19_15[5]\, N_1047_25, 
        \state_ns_i_a2_0_a4_0_19_12[5]\, 
        \state_ns_i_a2_0_a4_0_19_11[5]\, N_1047_5, 
        \state_ns_i_a2_0_a4_0_25_4[5]\, 
        \state_ns_i_a2_0_a4_0_25_2[5]\, 
        \state_ns_i_a2_0_a4_0_25_1[5]\, 
        \state_ns_i_a2_0_a4_0_25_0[5]\, 
        count_send_time_e2_0_a2_0_0, un1_state_13_0_a4_0_0, 
        \state[1]_net_1\, \state[3]_net_1\, 
        \state_ns_i_a2_0_a4_0_19_9_0[5]\, 
        \count_send_time_RNO[14]_net_1\, 
        \count_send_time_RNO[15]_net_1\, N_1092, 
        \count_send_time_RNO[16]_net_1\, 
        \count_send_time_RNO[6]_net_1\, N_1253, N_1230, 
        \count_send_time_RNO[7]_net_1\, \state_ns[6]\, 
        count_send_time_e10, N_1270, N_1272, N_1273, 
        count_send_time_e9, N_1265, N_1267, N_1268, 
        count_send_time_e8, N_1260, N_1262, N_1263, 
        count_send_time_e3, N_1249, N_1247, N_1246, 
        count_send_time_e2, N_1244, N_1242, N_1241, 
        count_send_time_e1, N_1239, N_1237, N_1236, 
        count_send_time_e11, N_1167, N_1169, N_1170, 
        count_send_time_e13, N_1086, N_1085, N_1087, 
        count_send_time_e12, N_1081, N_1080, N_1082, 
        \state_RNO[6]_net_1\, N_1027, N_1036, N_812, 
        \state[0]_net_1\, N_1037, un5_time_write, 
        \sel_data[1]_net_1\, \un13_time_write\, \un20_time_write\, 
        un27_time_write, un7_time_write, \time_write\, 
        un15_time_write, un22_time_write, un29_time_write, 
        un2_status_full_ack, un7_status_full_ack, 
        un12_status_full_ack, un17_status_full_ack, \data_ren\, 
        N_200, N_249, \time_select\, \time_ren\, 
        \update_and_sel_1[6]\, \update[0]_net_1\, 
        \update_and_sel_1[7]\, \update[1]_net_1\, 
        \update_and_sel_3[4]\, \update_and_sel_3[5]\, 
        \update_and_sel_5[2]\, \update_and_sel_5[3]\, 
        \update_and_sel_7[0]\, \update_and_sel_7[1]\, 
        \data_address[0]\, N_1279, N_1297, \data_address[1]\, 
        N_1280, N_1298, \data_address[2]\, N_1323, N_1299, 
        \data_address[3]\, N_1324, N_1300, \data_address[4]\, 
        N_1325, N_1301, \data_address[5]\, N_1326, N_1288, 
        \data_address[6]\, N_1327, N_1289, \data_address[7]\, 
        N_1328, N_1290, \data_address[8]\, N_1329, N_1291, 
        \data_address[9]\, N_1316, N_1292, \data_address[10]\, 
        N_1317, N_1293, \data_address[11]\, N_1318, N_1294, 
        \data_address[12]\, N_1319, N_1281, \data_address[13]\, 
        N_1320, N_1282, \data_address[14]\, N_1321, N_1283, 
        \sel_data[0]_net_1\, \data_address[15]\, N_1322, N_1284, 
        \data_address[16]\, N_1309, N_1285, \data_address[17]\, 
        N_1310, N_1286, \data_address[18]\, N_1311, N_1287, 
        \data_address[19]\, N_1312, N_902, \data_address[20]\, 
        N_1313, N_903, \data_address[21]\, N_1314, N_904, 
        \data_address[22]\, N_1315, N_905, \data_address[23]\, 
        N_1302, N_906, \data_address[24]\, N_1303, N_907, 
        \data_address[25]\, N_1304, N_908, \data_address[26]\, 
        N_1305, N_909, \data_address[27]\, N_1306, N_910, 
        \data_address[28]\, N_1307, N_911, \data_address[29]\, 
        N_1308, N_912, \data_address[30]\, N_1295, N_913, 
        \data_address[31]\, N_1296, N_914, N_1024, 
        \time_already_send[3]\, \time_already_send[2]\, N_1025, 
        \time_already_send[1]\, \count_send_time_RNO_1[6]_net_1\, 
        count_send_time_e0, \count_send_time_RNO[4]_net_1\, 
        N_1227, \count_send_time_RNO[5]_net_1\, N_1228, 
        \state_RNO_1[0]\, un1_data_send_ok, N_815, N_1040, N_1014, 
        \state_RNO[7]_net_1\, \time_fifo_ren\, N_1030, 
        un1_state_12, \state[6]_net_1\, \time_already_send[0]\, 
        \state_RNO_2[3]\, N_1033, \state_RNO_0[4]_net_1\, N_1044, 
        \state_RNO[5]_net_1\, N_1042, un1_state_13, 
        un1_time_send_ok, \state[5]_net_1\, time_send_0_sqmuxa, 
        update_0_sqmuxa, \time_send\, \data_send\, 
        \send_16_3_time[2]_net_1\, \send_16_3_time[1]_net_1\, 
        \un7_dmain[66]\, Ready, N_1012, Grant, OKAY, Fault, 
        N_1011, N_1013, N_960, N_959, N_958, N_957, N_964, N_963, 
        N_962, N_961, N_955, N_954, N_953, N_952, N_951, N_950, 
        N_949, N_948, N_947, N_956, N_965, N_966, N_967, N_968, 
        N_969, N_970, N_971, N_972, N_973, N_974, N_975, N_976, 
        N_977, N_978, Lock, Request, Store, 
        \addr_data_vector[97]\, \addr_data_vector[96]\, 
        \addr_data_vector[63]\, \addr_data_vector[61]\, 
        \addr_data_vector[60]\, \addr_data_vector[58]\, 
        \addr_data_vector[56]\, \addr_data_vector[36]\, 
        \addr_data_vector[42]\, \addr_data_vector[40]\, 
        \addr_data_vector[39]\, \addr_data_vector[38]\, 
        \addr_data_vector[37]\, \addr_data_vector[50]\, 
        \addr_data_vector[48]\, \addr_data_vector[46]\, 
        \addr_data_vector[44]\, \addr_data_vector[99]\, 
        \addr_data_vector[126]\, \addr_data_vector[123]\, 
        \addr_data_vector[121]\, \addr_data_vector[98]\, 
        \addr_data_vector[105]\, \addr_data_vector[109]\, 
        \addr_data_vector[107]\, \addr_data_vector[113]\, 
        \addr_data_vector[115]\, \addr_data_vector[118]\, 
        \addr_data_vector[119]\, \addr_data_vector[111]\, 
        \addr_data_vector[116]\, \addr_data_vector[117]\, 
        \addr_data_vector[65]\, \addr_data_vector[64]\, 
        \addr_data_vector[8]\, \addr_data_vector[7]\, 
        \addr_data_vector[6]\, \addr_data_vector[3]\, 
        \addr_data_vector[15]\, \addr_data_vector[14]\, 
        \addr_data_vector[12]\, \addr_data_vector[10]\, 
        \addr_data_vector[9]\, \addr_data_vector[29]\, 
        \addr_data_vector[27]\, \addr_data_vector[25]\, 
        \addr_data_vector[31]\, \addr_data_vector[69]\, 
        \addr_data_vector[68]\, \addr_data_vector[94]\, 
        \addr_data_vector[92]\, \addr_data_vector[90]\, 
        \addr_data_vector[66]\, \addr_data_vector[75]\, 
        \addr_data_vector[77]\, \addr_data_vector[82]\, 
        \addr_data_vector[81]\, \addr_data_vector[84]\, 
        \addr_data_vector[83]\, \addr_data_vector[87]\, 
        \addr_data_vector[88]\, \addr_data_vector[80]\, 
        \addr_data_vector[85]\, \addr_data_vector[86]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

    for all : \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\
	Use entity work.
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\(DEF_ARCH);
    for all : \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\
	Use entity work.
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\(DEF_ARCH);
    for all : lpp_dma_send_16word
	Use entity work.lpp_dma_send_16word(DEF_ARCH);
    for all : \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\
	Use entity work.
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\(DEF_ARCH);
    for all : lpp_dma_send_1word
	Use entity work.lpp_dma_send_1word(DEF_ARCH);
    for all : \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\
	Use entity work.
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\(DEF_ARCH);
    for all : DMA2AHB
	Use entity work.DMA2AHB(DEF_ARCH);
begin 

    time_ren_1z <= \time_ren\;
    data_ren_1z <= \data_ren\;
    un20_time_write <= \un20_time_write\;
    un13_time_write <= \un13_time_write\;

    \state[0]\ : DFN1C0
      port map(D => \state_RNO_1[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[0]_net_1\);
    
    \count_send_time_RNO_0[9]\ : OR3C
      port map(A => \state_0[2]_net_1\, B => 
        \count_send_time[9]_net_1\, C => N_1225, Y => N_1265);
    
    \count_send_time_RNO_4[30]\ : OR3C
      port map(A => N_1075, B => \count_send_time[30]_net_1\, C
         => N_1091, Y => N_1125);
    
    \sel_data[0]\ : DFN1E1C0
      port map(D => N_1016_i_0, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \state[7]_net_1\, Q => \sel_data[0]_net_1\);
    
    \gen_select_address.2.lpp_waveform_dma_selectaddress_I\ : 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_1\
      port map(nb_burst_available(10) => nb_burst_available(10), 
        nb_burst_available(9) => nb_burst_available(9), 
        nb_burst_available(8) => nb_burst_available(8), 
        nb_burst_available(7) => nb_burst_available(7), 
        nb_burst_available(6) => nb_burst_available(6), 
        nb_burst_available(5) => nb_burst_available(5), 
        nb_burst_available(4) => nb_burst_available(4), 
        nb_burst_available(3) => nb_burst_available(3), 
        nb_burst_available(2) => nb_burst_available(2), 
        nb_burst_available(1) => nb_burst_available(1), 
        nb_burst_available(0) => nb_burst_available(0), 
        status_full_err(2) => status_full_err(2), status_full(2)
         => status_full(2), sel_data(1) => \sel_data[1]_net_1\, 
        sel_data_1(1) => \sel_data_1[1]_net_1\, sel_data_0(1) => 
        \sel_data_0[1]_net_1\, update_and_sel_3(5) => 
        \update_and_sel_3[5]\, update_and_sel_3(4) => 
        \update_and_sel_3[4]\, addr_data_f2(31) => 
        addr_data_f2(31), addr_data_f2(30) => addr_data_f2(30), 
        addr_data_f2(29) => addr_data_f2(29), addr_data_f2(28)
         => addr_data_f2(28), addr_data_f2(27) => 
        addr_data_f2(27), addr_data_f2(26) => addr_data_f2(26), 
        addr_data_f2(25) => addr_data_f2(25), addr_data_f2(24)
         => addr_data_f2(24), addr_data_f2(23) => 
        addr_data_f2(23), addr_data_f2(22) => addr_data_f2(22), 
        addr_data_f2(21) => addr_data_f2(21), addr_data_f2(20)
         => addr_data_f2(20), addr_data_f2(19) => 
        addr_data_f2(19), addr_data_f2(18) => addr_data_f2(18), 
        addr_data_f2(17) => addr_data_f2(17), addr_data_f2(16)
         => addr_data_f2(16), addr_data_f2(15) => 
        addr_data_f2(15), addr_data_f2(14) => addr_data_f2(14), 
        addr_data_f2(13) => addr_data_f2(13), addr_data_f2(12)
         => addr_data_f2(12), addr_data_f2(11) => 
        addr_data_f2(11), addr_data_f2(10) => addr_data_f2(10), 
        addr_data_f2(9) => addr_data_f2(9), addr_data_f2(8) => 
        addr_data_f2(8), addr_data_f2(7) => addr_data_f2(7), 
        addr_data_f2(6) => addr_data_f2(6), addr_data_f2(5) => 
        addr_data_f2(5), addr_data_f2(4) => addr_data_f2(4), 
        addr_data_f2(3) => addr_data_f2(3), addr_data_f2(2) => 
        addr_data_f2(2), addr_data_f2(1) => addr_data_f2(1), 
        addr_data_f2(0) => addr_data_f2(0), status_full_ack(2)
         => status_full_ack(2), addr_data_vector_62 => 
        \addr_data_vector[65]\, addr_data_vector_61 => 
        \addr_data_vector[64]\, addr_data_vector_5 => 
        \addr_data_vector[8]\, addr_data_vector_4 => 
        \addr_data_vector[7]\, addr_data_vector_3 => 
        \addr_data_vector[6]\, addr_data_vector_0 => 
        \addr_data_vector[3]\, addr_data_vector_12 => 
        \addr_data_vector[15]\, addr_data_vector_11 => 
        \addr_data_vector[14]\, addr_data_vector_9 => 
        \addr_data_vector[12]\, addr_data_vector_7 => 
        \addr_data_vector[10]\, addr_data_vector_6 => 
        \addr_data_vector[9]\, addr_data_vector_26 => 
        \addr_data_vector[29]\, addr_data_vector_24 => 
        \addr_data_vector[27]\, addr_data_vector_22 => 
        \addr_data_vector[25]\, addr_data_vector_28 => 
        \addr_data_vector[31]\, addr_data_vector_66 => 
        \addr_data_vector[69]\, addr_data_vector_65 => 
        \addr_data_vector[68]\, addr_data_vector_91 => 
        \addr_data_vector[94]\, addr_data_vector_89 => 
        \addr_data_vector[92]\, addr_data_vector_87 => 
        \addr_data_vector[90]\, addr_data_vector_63 => 
        \addr_data_vector[66]\, addr_data_vector_72 => 
        \addr_data_vector[75]\, addr_data_vector_74 => 
        \addr_data_vector[77]\, addr_data_vector_79 => 
        \addr_data_vector[82]\, addr_data_vector_78 => 
        \addr_data_vector[81]\, addr_data_vector_81 => 
        \addr_data_vector[84]\, addr_data_vector_80 => 
        \addr_data_vector[83]\, addr_data_vector_84 => 
        \addr_data_vector[87]\, addr_data_vector_85 => 
        \addr_data_vector[88]\, addr_data_vector_77 => 
        \addr_data_vector[80]\, addr_data_vector_82 => 
        \addr_data_vector[85]\, addr_data_vector_83 => 
        \addr_data_vector[86]\, N_1329 => N_1329, N_1328 => 
        N_1328, N_1327 => N_1327, N_1324 => N_1324, N_1322 => 
        N_1322, N_1321 => N_1321, N_1319 => N_1319, N_1317 => 
        N_1317, N_1316 => N_1316, N_1308 => N_1308, N_1306 => 
        N_1306, N_1304 => N_1304, N_1296 => N_1296, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    \count_send_time_RNIRUBI[20]\ : NOR3C
      port map(A => count_send_time_e25_0_o3_m6_0_a2_2, B => 
        count_send_time_e25_0_o3_m6_0_a2_1, C => 
        count_send_time_e25_0_o3_m6_0_a2_6, Y => 
        count_send_time_e25_0_o3_m6_0_a2_7);
    
    \count_send_time_RNO_0[16]\ : OAI1
      port map(A => N_1077, B => \count_send_time[16]_net_1\, C
         => N_1091, Y => count_send_time_e16_i_0);
    
    \count_send_time_RNO_2[1]\ : OR2B
      port map(A => \count_send_time[1]_net_1\, B => N_1220, Y
         => N_1236);
    
    \count_send_time_RNO[4]\ : XA1A
      port map(A => N_1227, B => \count_send_time[4]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[4]_net_1\);
    
    \count_send_time_RNINOP61[10]\ : OR3B
      port map(A => \count_send_time[9]_net_1\, B => 
        \count_send_time[10]_net_1\, C => N_1225, Y => N_1159);
    
    \gen_select_address.0.lpp_waveform_dma_selectaddress_I\ : 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_3\
      port map(nb_burst_available(10) => nb_burst_available(10), 
        nb_burst_available(9) => nb_burst_available(9), 
        nb_burst_available(8) => nb_burst_available(8), 
        nb_burst_available(7) => nb_burst_available(7), 
        nb_burst_available(6) => nb_burst_available(6), 
        nb_burst_available(5) => nb_burst_available(5), 
        nb_burst_available(4) => nb_burst_available(4), 
        nb_burst_available(3) => nb_burst_available(3), 
        nb_burst_available(2) => nb_burst_available(2), 
        nb_burst_available(1) => nb_burst_available(1), 
        nb_burst_available(0) => nb_burst_available(0), 
        status_full_err(0) => status_full_err(0), status_full(0)
         => status_full(0), sel_data(1) => \sel_data[1]_net_1\, 
        sel_data_1(1) => \sel_data_1[1]_net_1\, sel_data_0(1) => 
        \sel_data_0[1]_net_1\, update_and_sel_7(1) => 
        \update_and_sel_7[1]\, update_and_sel_7(0) => 
        \update_and_sel_7[0]\, addr_data_f0(31) => 
        addr_data_f0(31), addr_data_f0(30) => addr_data_f0(30), 
        addr_data_f0(29) => addr_data_f0(29), addr_data_f0(28)
         => addr_data_f0(28), addr_data_f0(27) => 
        addr_data_f0(27), addr_data_f0(26) => addr_data_f0(26), 
        addr_data_f0(25) => addr_data_f0(25), addr_data_f0(24)
         => addr_data_f0(24), addr_data_f0(23) => 
        addr_data_f0(23), addr_data_f0(22) => addr_data_f0(22), 
        addr_data_f0(21) => addr_data_f0(21), addr_data_f0(20)
         => addr_data_f0(20), addr_data_f0(19) => 
        addr_data_f0(19), addr_data_f0(18) => addr_data_f0(18), 
        addr_data_f0(17) => addr_data_f0(17), addr_data_f0(16)
         => addr_data_f0(16), addr_data_f0(15) => 
        addr_data_f0(15), addr_data_f0(14) => addr_data_f0(14), 
        addr_data_f0(13) => addr_data_f0(13), addr_data_f0(12)
         => addr_data_f0(12), addr_data_f0(11) => 
        addr_data_f0(11), addr_data_f0(10) => addr_data_f0(10), 
        addr_data_f0(9) => addr_data_f0(9), addr_data_f0(8) => 
        addr_data_f0(8), addr_data_f0(7) => addr_data_f0(7), 
        addr_data_f0(6) => addr_data_f0(6), addr_data_f0(5) => 
        addr_data_f0(5), addr_data_f0(4) => addr_data_f0(4), 
        addr_data_f0(3) => addr_data_f0(3), addr_data_f0(2) => 
        addr_data_f0(2), addr_data_f0(1) => addr_data_f0(1), 
        addr_data_f0(0) => addr_data_f0(0), status_full_ack(0)
         => status_full_ack(0), addr_data_vector_69 => 
        \addr_data_vector[69]\, addr_data_vector_68 => 
        \addr_data_vector[68]\, addr_data_vector_66 => 
        \addr_data_vector[66]\, addr_data_vector_77 => 
        \addr_data_vector[77]\, addr_data_vector_75 => 
        \addr_data_vector[75]\, addr_data_vector_86 => 
        \addr_data_vector[86]\, addr_data_vector_85 => 
        \addr_data_vector[85]\, addr_data_vector_84 => 
        \addr_data_vector[84]\, addr_data_vector_83 => 
        \addr_data_vector[83]\, addr_data_vector_82 => 
        \addr_data_vector[82]\, addr_data_vector_81 => 
        \addr_data_vector[81]\, addr_data_vector_80 => 
        \addr_data_vector[80]\, addr_data_vector_92 => 
        \addr_data_vector[92]\, addr_data_vector_90 => 
        \addr_data_vector[90]\, addr_data_vector_88 => 
        \addr_data_vector[88]\, addr_data_vector_87 => 
        \addr_data_vector[87]\, addr_data_vector_94 => 
        \addr_data_vector[94]\, addr_data_vector_65 => 
        \addr_data_vector[65]\, addr_data_vector_64 => 
        \addr_data_vector[64]\, addr_data_vector_3 => 
        \addr_data_vector[3]\, addr_data_vector_31 => 
        \addr_data_vector[31]\, addr_data_vector_14 => 
        \addr_data_vector[14]\, addr_data_vector_15 => 
        \addr_data_vector[15]\, addr_data_vector_27 => 
        \addr_data_vector[27]\, addr_data_vector_29 => 
        \addr_data_vector[29]\, addr_data_vector_25 => 
        \addr_data_vector[25]\, addr_data_vector_6 => 
        \addr_data_vector[6]\, addr_data_vector_8 => 
        \addr_data_vector[8]\, addr_data_vector_7 => 
        \addr_data_vector[7]\, addr_data_vector_10 => 
        \addr_data_vector[10]\, addr_data_vector_9 => 
        \addr_data_vector[9]\, addr_data_vector_12 => 
        \addr_data_vector[12]\, N_1326 => N_1326, N_1325 => 
        N_1325, N_1323 => N_1323, N_1320 => N_1320, N_1318 => 
        N_1318, N_1315 => N_1315, N_1314 => N_1314, N_1313 => 
        N_1313, N_1312 => N_1312, N_1311 => N_1311, N_1310 => 
        N_1310, N_1309 => N_1309, N_1307 => N_1307, N_1305 => 
        N_1305, N_1303 => N_1303, N_1302 => N_1302, N_1295 => 
        N_1295, N_1280 => N_1280, N_1279 => N_1279, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    \count_send_time_RNIFF6R1[20]\ : OR3C
      port map(A => N_1063, B => \count_send_time[19]_net_1\, C
         => \count_send_time[20]_net_1\, Y => N_1066);
    
    \sel_data_0_RNI0MA8[0]\ : OR2B
      port map(A => \sel_data[1]_net_1\, B => 
        \sel_data_0[0]_net_1\, Y => un5_time_write);
    
    \count_send_time_RNO[26]\ : XA1A
      port map(A => N_1163, B => \count_send_time[26]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[26]_net_1\);
    
    \count_send_time_RNINK24[24]\ : NOR2B
      port map(A => \count_send_time[24]_net_1\, B => 
        \count_send_time[18]_net_1\, Y => 
        count_send_time_e25_0_o3_m6_0_a2_1);
    
    \sel_data_RNIM70E[0]\ : MX2C
      port map(A => N_1308, B => N_912, S => \sel_data[0]_net_1\, 
        Y => \data_address[29]\);
    
    \all_time_write.0.time_already_send_RNI944DP[0]\ : MX2
      port map(A => N_1025, B => \time_already_send[0]\, S => 
        ready_i_0(0), Y => N_1026);
    
    \count_send_time[0]\ : DFN1
      port map(D => count_send_time_e0, CLK => HCLK_c, Q => 
        \count_send_time[0]_net_1\);
    
    \count_send_time_RNO_3[2]\ : OR3B
      port map(A => \count_send_time[0]_net_1\, B => 
        \count_send_time[1]_net_1\, C => 
        \count_send_time[2]_net_1\, Y => 
        count_send_time_e2_0_a2_1_0);
    
    \count_send_time_RNO_0[10]\ : AO1C
      port map(A => N_1225, B => \count_send_time[9]_net_1\, C
         => count_send_time_e10_0_a2_0, Y => N_1270);
    
    \count_send_time_RNO[2]\ : OR3C
      port map(A => N_1244, B => N_1242, C => N_1241, Y => 
        count_send_time_e2);
    
    time_fifo_ren_RNO : INV
      port map(A => time_fifo_ren_1, Y => time_fifo_ren_1_i);
    
    lpp_dma_send_16word_1 : lpp_dma_send_16word
      port map(un7_dmain(66) => \un7_dmain[66]\, data_address(31)
         => \data_address[31]\, data_address(30) => 
        \data_address[30]\, data_address(29) => 
        \data_address[29]\, data_address(28) => 
        \data_address[28]\, data_address(27) => 
        \data_address[27]\, data_address(26) => 
        \data_address[26]\, data_address(25) => 
        \data_address[25]\, data_address(24) => 
        \data_address[24]\, data_address(23) => 
        \data_address[23]\, data_address(22) => 
        \data_address[22]\, data_address(21) => 
        \data_address[21]\, data_address(20) => 
        \data_address[20]\, data_address(19) => 
        \data_address[19]\, data_address(18) => 
        \data_address[18]\, data_address(17) => 
        \data_address[17]\, data_address(16) => 
        \data_address[16]\, data_address(15) => 
        \data_address[15]\, data_address(14) => 
        \data_address[14]\, data_address(13) => 
        \data_address[13]\, data_address(12) => 
        \data_address[12]\, data_address(11) => 
        \data_address[11]\, data_address(10) => 
        \data_address[10]\, data_address(9) => \data_address[9]\, 
        data_address(8) => \data_address[8]\, data_address(7) => 
        \data_address[7]\, data_address(6) => \data_address[6]\, 
        data_address(5) => \data_address[5]\, data_address(4) => 
        \data_address[4]\, data_address(3) => \data_address[3]\, 
        data_address(2) => \data_address[2]\, data_address(1) => 
        \data_address[1]\, data_address(0) => \data_address[0]\, 
        Store => Store, Fault => Fault, un1_data_send_ok => 
        un1_data_send_ok, Request_0 => Request, N_1011 => N_1011, 
        Lock_0 => Lock, N_1013 => N_1013, N_957 => N_957, N_956
         => N_956, N_955 => N_955, N_954 => N_954, N_953 => N_953, 
        N_952 => N_952, N_951 => N_951, N_964 => N_964, N_963 => 
        N_963, N_962 => N_962, N_961 => N_961, N_960 => N_960, 
        time_select => \time_select\, N_959 => N_959, N_958 => 
        N_958, N_971 => N_971, N_970 => N_970, N_969 => N_969, 
        N_968 => N_968, N_967 => N_967, N_966 => N_966, N_965 => 
        N_965, N_978 => N_978, N_977 => N_977, N_976 => N_976, 
        N_975 => N_975, N_974 => N_974, N_973 => N_973, N_972 => 
        N_972, N_950 => N_950, N_949 => N_949, N_948 => N_948, 
        time_select_0 => \time_select_0\, N_947 => N_947, N_249
         => N_249, Grant => Grant, Ready => Ready, data_send => 
        \data_send\, OKAY => OKAY, N_200 => N_200, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    \count_send_time_RNO_1[6]\ : NOR3B
      port map(A => N_1219, B => \count_send_time[5]_net_1\, C
         => N_1145, Y => \count_send_time_RNO_1[6]_net_1\);
    
    \count_send_time_RNO_0[27]\ : OR2A
      port map(A => N_1146, B => N_1145, Y => N_1164);
    
    \count_send_time_RNO_1[19]\ : OR2B
      port map(A => \count_send_time[19]_net_1\, B => N_1220, Y
         => N_1102);
    
    \count_send_time_RNIRQ3N1[17]\ : NOR3C
      port map(A => N_1061, B => \count_send_time[17]_net_1\, C
         => \count_send_time[18]_net_1\, Y => N_1063);
    
    \count_send_time[14]\ : DFN1
      port map(D => \count_send_time_RNO[14]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[14]_net_1\);
    
    \state[6]\ : DFN1C0
      port map(D => \state_RNO[6]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[6]_net_1\);
    
    \count_send_time_RNO_2[18]\ : NOR2B
      port map(A => \count_send_time[18]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e18_0_a2_0_0);
    
    \count_send_time[21]\ : DFN1
      port map(D => count_send_time_e21, CLK => HCLK_c, Q => 
        \count_send_time[21]_net_1\);
    
    \count_send_time_RNO[14]\ : OA1C
      port map(A => N_1059, B => N_1145_0, C => 
        count_send_time_e14_i_0, Y => 
        \count_send_time_RNO[14]_net_1\);
    
    \count_send_time[31]\ : DFN1
      port map(D => count_send_time_e31, CLK => HCLK_c, Q => 
        \count_send_time[31]_net_1\);
    
    \update_RNIPECD_0[1]\ : NOR2A
      port map(A => \update[1]_net_1\, B => \un20_time_write\, Y
         => \update_and_sel_5[3]\);
    
    \sel_data_RNIP45D[0]\ : MX2C
      port map(A => N_1321, B => N_1283, S => \sel_data[0]_net_1\, 
        Y => \data_address[14]\);
    
    \count_send_time_RNI8KVA[2]\ : OR3C
      port map(A => \count_send_time[0]_net_1\, B => 
        \count_send_time[1]_net_1\, C => 
        \count_send_time[2]_net_1\, Y => N_1217);
    
    \count_send_time_RNO[22]\ : OR3C
      port map(A => N_1117, B => N_1118, C => N_1119, Y => 
        count_send_time_e22);
    
    time_write_RNO : AO1D
      port map(A => un1_state_13_0_a4_0_0, B => \state[7]_net_1\, 
        C => N_1033, Y => un1_state_13);
    
    \count_send_time[17]\ : DFN1
      port map(D => \count_send_time_RNO[17]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[17]_net_1\);
    
    \state_RNIKSS3_0[2]\ : OAI1
      port map(A => \state[2]_net_1\, B => \state[7]_net_1\, C
         => HRESETn_c, Y => N_1220);
    
    \count_send_time_RNO_0[3]\ : OR3
      port map(A => N_1217, B => \count_send_time[3]_net_1\, C
         => N_1145_0, Y => N_1249);
    
    \all_data_ren.2.data_time_ren_3[2]\ : OR2A
      port map(A => \time_ren\, B => \un13_time_write\, Y => 
        time_ren(2));
    
    \all_data_ren.1.data_data_ren_5[1]\ : OR2A
      port map(A => \data_ren\, B => \un20_time_write\, Y => 
        data_ren(1));
    
    \count_send_time_RNO_2[8]\ : OR3B
      port map(A => N_1223, B => \count_send_time[7]_net_1\, C
         => count_send_time_e8_0_a2_1_0, Y => N_1263);
    
    \count_send_time_RNIN9B7[4]\ : NOR2
      port map(A => \count_send_time[4]_net_1\, B => 
        \count_send_time[5]_net_1\, Y => 
        \state_ns_i_a2_0_a4_0_25_0[5]\);
    
    \update_RNIOECD_1[0]\ : OR2A
      port map(A => \update[0]_net_1\, B => \un13_time_write\, Y
         => \update_and_sel_3[4]\);
    
    \state_ns_i_a2_0_a3_0[5]\ : NAND2
      port map(A => N_1026, B => \state[4]_net_1\, Y => N_1049);
    
    \sel_data_0_RNIKH5P[0]\ : MX2C
      port map(A => N_1324, B => N_1300, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[3]\);
    
    \count_send_time_RNO[7]\ : XA1
      port map(A => N_1230, B => \count_send_time[7]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[7]_net_1\);
    
    \count_send_time_RNO_2[9]\ : OR3
      port map(A => N_1145_0, B => \count_send_time[9]_net_1\, C
         => N_1225, Y => N_1268);
    
    \sel_data_0_RNIKIAC[0]\ : MX2C
      port map(A => N_1319, B => N_1281, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[12]\);
    
    \count_send_time[25]\ : DFN1
      port map(D => count_send_time_e25, CLK => HCLK_c, Q => 
        \count_send_time[25]_net_1\);
    
    \update_RNIPECD[1]\ : NOR2A
      port map(A => \update[1]_net_1\, B => un5_time_write, Y => 
        \update_and_sel_1[7]\);
    
    \count_send_time[5]\ : DFN1
      port map(D => \count_send_time_RNO[5]_net_1\, CLK => HCLK_c, 
        Q => \count_send_time[5]_net_1\);
    
    \update[1]\ : DFN1E0C0
      port map(D => \state[0]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_12, Q => \update[1]_net_1\);
    
    time_select : DFN1E1C0
      port map(D => time_fifo_ren_1, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_816, Q => \time_select\);
    
    \count_send_time_RNO_0[2]\ : OR2
      port map(A => count_send_time_e2_0_a2_1_0, B => N_1145_0, Y
         => N_1244);
    
    \count_send_time_RNO[27]\ : XA1A
      port map(A => N_1164, B => \count_send_time[27]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[27]_net_1\);
    
    \update_RNIOECD_0[0]\ : OR2A
      port map(A => \update[0]_net_1\, B => \un20_time_write\, Y
         => \update_and_sel_5[2]\);
    
    \state_RNIHU8A[3]\ : NOR2A
      port map(A => \state[3]_net_1\, B => un1_time_send_ok, Y
         => N_1033);
    
    \sel_data_RNIU60E[0]\ : MX2C
      port map(A => N_1302, B => N_906, S => \sel_data[0]_net_1\, 
        Y => \data_address[23]\);
    
    \count_send_time_RNO_1[10]\ : OR2B
      port map(A => \count_send_time[10]_net_1\, B => N_1220, Y
         => N_1272);
    
    \count_send_time_RNO[0]\ : MX2A
      port map(A => N_1145, B => N_1220, S => 
        \count_send_time[0]_net_1\, Y => count_send_time_e0);
    
    \count_send_time_RNO[10]\ : OR3C
      port map(A => N_1270, B => N_1272, C => N_1273, Y => 
        count_send_time_e10);
    
    \all_time_write.3.time_already_send[3]\ : DFN1E1C0
      port map(D => un7_time_write, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un2_status_full_ack, Q => 
        \time_already_send[3]\);
    
    \sel_data_0[1]\ : DFN1E1C0
      port map(D => N_1015, CLK => HCLK_c, CLR => HRESETn_c, E
         => \state[7]_net_1\, Q => \sel_data_0[1]_net_1\);
    
    \count_send_time_RNO_4[12]\ : OR2
      port map(A => \count_send_time[12]_net_1\, B => N_1145_0, Y
         => count_send_time_e12_0_a2_1_0);
    
    \count_send_time_RNI4A1J1[16]\ : NOR3C
      port map(A => N_1059, B => \count_send_time[15]_net_1\, C
         => \count_send_time[16]_net_1\, Y => N_1061);
    
    \state[4]\ : DFN1C0
      port map(D => \state_RNO_0[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \state[4]_net_1\);
    
    time_write : DFN1E0C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_13, Q => \time_write\);
    
    data_send_RNO : NOR3
      port map(A => \state[0]_net_1\, B => \state[1]_net_1\, C
         => \state[7]_net_1\, Y => N_812);
    
    \sel_data_1[1]\ : DFN1E1C0
      port map(D => N_1015, CLK => HCLK_c, CLR => HRESETn_c, E
         => \state[7]_net_1\, Q => \sel_data_1[1]_net_1\);
    
    \sel_data_0_RNIBH4P[0]\ : MX2C
      port map(A => N_1280, B => N_1298, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[1]\);
    
    \count_send_time[28]\ : DFN1
      port map(D => \count_send_time_RNO[28]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[28]_net_1\);
    
    \update_RNIOECD[0]\ : OR2A
      port map(A => \update[0]_net_1\, B => un5_time_write, Y => 
        \update_and_sel_1[6]\);
    
    \sel_data_RNIANVD[0]\ : MX2C
      port map(A => N_1312, B => N_902, S => \sel_data[0]_net_1\, 
        Y => \data_address[19]\);
    
    \count_send_time_RNIGL6A[22]\ : NOR3C
      port map(A => \count_send_time[22]_net_1\, B => 
        \count_send_time[21]_net_1\, C => 
        count_send_time_e25_0_o3_m6_0_a2_4, Y => 
        count_send_time_e25_0_o3_m6_0_a2_6);
    
    \count_send_time[8]\ : DFN1
      port map(D => count_send_time_e8, CLK => HCLK_c, Q => 
        \count_send_time[8]_net_1\);
    
    \sel_data_0_RNIO31Q[0]\ : MX2C
      port map(A => N_1326, B => N_1288, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[5]\);
    
    \count_send_time_RNO[13]\ : OR3C
      port map(A => N_1086, B => N_1085, C => N_1087, Y => 
        count_send_time_e13);
    
    \state[7]\ : DFN1P0
      port map(D => \state_RNO[7]_net_1\, CLK => HCLK_c, PRE => 
        HRESETn_c, Q => \state[7]_net_1\);
    
    \count_send_time_RNIT09T[6]\ : NOR2A
      port map(A => N_1223, B => N_1145, Y => N_1230);
    
    \count_send_time_RNO[3]\ : OR3C
      port map(A => N_1249, B => N_1247, C => N_1246, Y => 
        count_send_time_e3);
    
    \count_send_time[10]\ : DFN1
      port map(D => count_send_time_e10, CLK => HCLK_c, Q => 
        \count_send_time[10]_net_1\);
    
    time_write_RNI6IL9_2 : NOR2A
      port map(A => \time_write\, B => un27_time_write, Y => 
        un29_time_write);
    
    \count_send_time_RNO_2[30]\ : OR3B
      port map(A => N_1146, B => \count_send_time[27]_net_1\, C
         => count_send_time_e30_0_a2_2_1, Y => N_1128);
    
    \state[5]\ : DFN1C0
      port map(D => \state_RNO[5]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[5]_net_1\);
    
    data_send : DFN1E0C0
      port map(D => \state[1]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_812, Q => \data_send\);
    
    \count_send_time_RNI9946[30]\ : OR2A
      port map(A => \count_send_time[30]_net_1\, B => N_1075, Y
         => N_1161);
    
    \DMAWriteFSM_p.sel_data_3_i_a4[0]\ : OR2A
      port map(A => ready_i_0(2), B => ready_i_0(1), Y => N_1037);
    
    \sel_data_0_RNIG15P[0]\ : MX2C
      port map(A => N_1323, B => N_1299, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[2]\);
    
    \update_RNIPECD_2[1]\ : NOR2A
      port map(A => \update[1]_net_1\, B => un27_time_write, Y
         => \update_and_sel_7[1]\);
    
    \count_send_time_RNO_1[2]\ : OR2B
      port map(A => count_send_time_e2_0_a2_0_0, B => 
        \state_0[2]_net_1\, Y => N_1242);
    
    \state_RNIMMJ[4]\ : NOR2
      port map(A => \state[6]_net_1\, B => \state[4]_net_1\, Y
         => N_1030);
    
    GND_i : GND
      port map(Y => \GND\);
    
    time_send_RNO : NOR2
      port map(A => N_1030, B => N_1026, Y => time_send_0_sqmuxa);
    
    \sel_data_0_RNI0MA8_1[0]\ : OR2A
      port map(A => \sel_data[1]_net_1\, B => 
        \sel_data_0[0]_net_1\, Y => \un13_time_write\);
    
    \count_send_time_RNO_3[24]\ : NOR2B
      port map(A => \count_send_time[24]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e24_0_a2_0_0);
    
    \count_send_time_RNO_0[25]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[25]_net_1\, C => 
        count_send_time_e25_0_o3_N_7_i_0, Y => N_1178);
    
    \count_send_time_RNO_3[12]\ : NOR2B
      port map(A => \count_send_time[12]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e12_0_a2_0_0);
    
    \count_send_time_RNIRPB7[6]\ : NOR2
      port map(A => \count_send_time[6]_net_1\, B => 
        \count_send_time[7]_net_1\, Y => 
        \state_ns_i_a2_0_a4_0_25_1[5]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \DMAWriteFSM_p.sel_data_3_i[0]\ : NOR3B
      port map(A => N_1037, B => N_1027, C => ready_i_0(0), Y => 
        N_1016_i_0);
    
    \state_RNO_0[5]\ : OR2A
      port map(A => \state[5]_net_1\, B => un1_time_send_ok, Y
         => N_1042);
    
    \state_RNO_0[4]\ : OR2B
      port map(A => \state[5]_net_1\, B => un1_time_send_ok, Y
         => N_1044);
    
    \sel_data_RNITM0E[0]\ : MX2C
      port map(A => N_1295, B => N_913, S => \sel_data[0]_net_1\, 
        Y => \data_address[30]\);
    
    \count_send_time_RNO_3[31]\ : OR3B
      port map(A => N_1146, B => \count_send_time[27]_net_1\, C
         => N_1161, Y => N_1162);
    
    \sel_data_RNII70E[0]\ : MX2C
      port map(A => N_1307, B => N_911, S => \sel_data[0]_net_1\, 
        Y => \data_address[28]\);
    
    \count_send_time_RNO_1[25]\ : OR2B
      port map(A => \count_send_time[25]_net_1\, B => N_1220, Y
         => N_1177);
    
    \count_send_time_RNO_2[25]\ : OR3
      port map(A => N_1145_0, B => \count_send_time[25]_net_1\, C
         => count_send_time_e25_0_o3_N_7_i_0, Y => N_1180);
    
    \count_send_time_RNINO24[24]\ : OR2
      port map(A => \count_send_time[24]_net_1\, B => 
        \count_send_time[25]_net_1\, Y => state_tr13_0_a2_17_1);
    
    \DMAWriteFSM_p.sel_data_3_i_o3[0]\ : OR2A
      port map(A => ready_i_0(3), B => ready_i_0(1), Y => N_1027);
    
    \state_RNO_0[7]\ : OR3B
      port map(A => \send_16_3_time_1_sqmuxa_i_o3_0\, B => 
        \state[7]_net_1\, C => N_1027, Y => N_1040);
    
    \count_send_time[7]\ : DFN1
      port map(D => \count_send_time_RNO[7]_net_1\, CLK => HCLK_c, 
        Q => \count_send_time[7]_net_1\);
    
    \count_send_time_RNO[25]\ : OR3C
      port map(A => N_1178, B => N_1177, C => N_1180, Y => 
        count_send_time_e25);
    
    \count_send_time_RNO_1[9]\ : OR2B
      port map(A => \count_send_time[9]_net_1\, B => N_1220, Y
         => N_1267);
    
    \count_send_time_RNIVS36[16]\ : NOR3C
      port map(A => \count_send_time[17]_net_1\, B => 
        \count_send_time[16]_net_1\, C => 
        \count_send_time[23]_net_1\, Y => 
        count_send_time_e25_0_o3_m6_0_a2_4);
    
    \count_send_time_RNO[31]\ : OR3C
      port map(A => N_1191, B => N_1193, C => N_1194, Y => 
        count_send_time_e31);
    
    \state_ns_i_a2_0_RNO_2[5]\ : NOR2A
      port map(A => \state[7]_net_1\, B => 
        \send_16_3_time[0]_net_1\, Y => 
        \state_ns_i_a2_0_a3_0[5]_net_1\);
    
    \count_send_time_RNIM7MP[6]\ : NOR3C
      port map(A => N_1219, B => \count_send_time[5]_net_1\, C
         => \count_send_time[6]_net_1\, Y => N_1223);
    
    \state_RNO[1]\ : NOR3C
      port map(A => state_tr13_0_a2_14, B => N_1047_25, C => 
        state_tr13_0_a2_15, Y => \state_ns[6]\);
    
    \state_RNIKSS3[2]\ : OR3B
      port map(A => \state[7]_net_1\, B => HRESETn_c, C => 
        \state[2]_net_1\, Y => N_1091);
    
    \count_send_time_RNO_3[22]\ : NOR2B
      port map(A => \count_send_time[22]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e22_0_a2_0);
    
    \count_send_time_RNI6158[16]\ : OR3A
      port map(A => \state_ns_i_a2_0_a4_0_19_9_0[5]\, B => 
        \count_send_time[17]_net_1\, C => 
        \count_send_time[16]_net_1\, Y => state_tr13_0_a2_9);
    
    \count_send_time_RNO_0[13]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[13]_net_1\, C => N_1057, Y => N_1086);
    
    time_write_RNI6IL9 : NOR2A
      port map(A => \time_write\, B => un5_time_write, Y => 
        un7_time_write);
    
    \sel_data_0[0]\ : DFN1E1C0
      port map(D => N_1016_i_0, CLK => HCLK_c, CLR => HRESETn_c, 
        E => \state[7]_net_1\, Q => \sel_data_0[0]_net_1\);
    
    \count_send_time_RNO_0[14]\ : OAI1
      port map(A => \count_send_time_RNO_1[14]_net_1\, B => 
        \count_send_time[14]_net_1\, C => N_1091, Y => 
        count_send_time_e14_i_0);
    
    \sel_data_0_RNIGHOH_0[0]\ : OR2A
      port map(A => \time_ren\, B => un5_time_write, Y => 
        time_ren(3));
    
    \count_send_time_RNO[8]\ : OR3C
      port map(A => N_1260, B => N_1262, C => N_1263, Y => 
        count_send_time_e8);
    
    \count_send_time[26]\ : DFN1
      port map(D => \count_send_time_RNO[26]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[26]_net_1\);
    
    \state_RNIQLS[5]\ : NOR3
      port map(A => \state[3]_net_1\, B => \state[5]_net_1\, C
         => \state[0]_net_1\, Y => N_816);
    
    \state_RNILNKV11[7]\ : AO1C
      port map(A => N_1027, B => \send_16_3_time_1_sqmuxa_i_o3_0\, 
        C => \state[7]_net_1\, Y => N_1014);
    
    \count_send_time_RNIU2FB[29]\ : NOR3
      port map(A => \count_send_time[29]_net_1\, B => 
        \count_send_time[28]_net_1\, C => N_1047_5, Y => 
        state_tr13_0_a2_7);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \count_send_time_RNI5L58[22]\ : NOR3A
      port map(A => state_tr13_0_a2_6, B => 
        \count_send_time[22]_net_1\, C => 
        \count_send_time[21]_net_1\, Y => state_tr13_0_a2_10);
    
    \sel_data[1]\ : DFN1E1C0
      port map(D => N_1015, CLK => HCLK_c, CLR => HRESETn_c, E
         => \state[7]_net_1\, Q => \sel_data[1]_net_1\);
    
    \count_send_time_RNIV9C7[8]\ : OR2
      port map(A => \count_send_time[9]_net_1\, B => 
        \count_send_time[8]_net_1\, Y => N_1047_5);
    
    \all_time_write.0.time_already_send[0]\ : DFN1E1C0
      port map(D => un29_time_write, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un17_status_full_ack, Q => 
        \time_already_send[0]\);
    
    \sel_data_0_RNI4K2Q[0]\ : MX2C
      port map(A => N_1329, B => N_1291, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[8]\);
    
    \count_send_time_RNIKS24[30]\ : NOR2
      port map(A => \count_send_time[23]_net_1\, B => 
        \count_send_time[30]_net_1\, Y => state_tr13_0_a2_6);
    
    \count_send_time_RNI29SA1[12]\ : OR3B
      port map(A => \count_send_time[11]_net_1\, B => 
        \count_send_time[12]_net_1\, C => N_1159, Y => N_1057);
    
    \sel_data_0_RNIIPAU1_0[0]\ : OR2A
      port map(A => \data_ren\, B => un5_time_write, Y => 
        data_ren(3));
    
    \count_send_time[29]\ : DFN1
      port map(D => \count_send_time_RNO[29]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[29]_net_1\);
    
    \send_16_3_time[1]\ : DFN1E0C0
      port map(D => \send_16_3_time[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => N_1014, Q => 
        \send_16_3_time[1]_net_1\);
    
    \sel_data_RNI670E[0]\ : MX2C
      port map(A => N_1304, B => N_908, S => \sel_data[0]_net_1\, 
        Y => \data_address[25]\);
    
    \state_RNO[4]\ : AO1B
      port map(A => \state[6]_net_1\, B => N_1026, C => N_1044, Y
         => \state_RNO_0[4]_net_1\);
    
    \count_send_time_RNO[19]\ : OR3C
      port map(A => N_1103, B => N_1102, C => N_1104, Y => 
        count_send_time_e19);
    
    send_16_3_time_1_sqmuxa_i_o3_0 : NOR2
      port map(A => ready_i_0(2), B => ready_i_0(0), Y => 
        \send_16_3_time_1_sqmuxa_i_o3_0\);
    
    \all_time_write.3.time_already_send_RNO[3]\ : OR2
      port map(A => status_full_ack(3), B => un7_time_write, Y
         => un2_status_full_ack);
    
    \state_ns_i_a2_0_RNO_3[5]\ : OR3C
      port map(A => \state_ns_i_a2_0_a4_0_19_12[5]\, B => 
        \state_ns_i_a2_0_a4_0_19_11[5]\, C => 
        \state_ns_i_a2_0_a4_0_19_15[5]\, Y => 
        \state_ns_i_a2_0_a4_0_19_i[5]\);
    
    \sel_data_RNIA70E[0]\ : MX2C
      port map(A => N_1305, B => N_909, S => \sel_data[0]_net_1\, 
        Y => \data_address[26]\);
    
    \count_send_time_RNO_1[30]\ : AOI1B
      port map(A => \count_send_time[30]_net_1\, B => N_1220, C
         => N_1125, Y => count_send_time_e30_0_0);
    
    \count_send_time[13]\ : DFN1
      port map(D => count_send_time_e13, CLK => HCLK_c, Q => 
        \count_send_time[13]_net_1\);
    
    \count_send_time[12]\ : DFN1
      port map(D => count_send_time_e12, CLK => HCLK_c, Q => 
        \count_send_time[12]_net_1\);
    
    \sel_data_0_RNI0MA8_0[0]\ : OR2A
      port map(A => \sel_data_0[0]_net_1\, B => 
        \sel_data[1]_net_1\, Y => \un20_time_write\);
    
    \DMAWriteFSM_p.sel_data_3_i[1]\ : NOR3
      port map(A => N_1036, B => ready_i_0(0), C => ready_i_0(1), 
        Y => N_1015);
    
    \count_send_time_RNO_0[12]\ : AO1C
      port map(A => N_1159, B => \count_send_time[11]_net_1\, C
         => count_send_time_e12_0_a2_0_0, Y => N_1081);
    
    \count_send_time_RNO[24]\ : OR3C
      port map(A => N_1173, B => N_1172, C => N_1175, Y => 
        count_send_time_e24);
    
    \count_send_time_RNO_2[3]\ : OR2B
      port map(A => \count_send_time[3]_net_1\, B => N_1220, Y
         => N_1246);
    
    \sel_data_0_RNIGIAC[0]\ : MX2C
      port map(A => N_1318, B => N_1294, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[11]\);
    
    \count_send_time_RNI23LE[0]\ : NOR3B
      port map(A => \count_send_time[1]_net_1\, B => 
        \state_ns_i_a2_0_a4_0_25_2[5]\, C => 
        \count_send_time[0]_net_1\, Y => 
        \state_ns_i_a2_0_a4_0_25_4[5]\);
    
    time_fifo_ren_RNIGRD9 : NOR2A
      port map(A => \time_select\, B => \time_fifo_ren\, Y => 
        \time_ren\);
    
    \count_send_time_RNO_0[30]\ : AO1B
      port map(A => \count_send_time[27]_net_1\, B => N_1146, C
         => count_send_time_e30_0_a2_0_0, Y => N_1126);
    
    \count_send_time_RNO_1[13]\ : OR2B
      port map(A => \count_send_time[13]_net_1\, B => N_1220, Y
         => N_1085);
    
    \count_send_time_RNO_2[19]\ : OR3A
      port map(A => N_1063, B => N_1145, C => 
        \count_send_time[19]_net_1\, Y => N_1104);
    
    \count_send_time_RNO_1[14]\ : NOR3A
      port map(A => \count_send_time[13]_net_1\, B => N_1057, C
         => N_1145, Y => \count_send_time_RNO_1[14]_net_1\);
    
    \count_send_time_RNO_0[6]\ : NOR2
      port map(A => \count_send_time[6]_net_1\, B => 
        \count_send_time_RNO_1[6]_net_1\, Y => N_1253);
    
    \count_send_time_RNO_0[11]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[11]_net_1\, C => N_1159, Y => N_1167);
    
    \count_send_time_RNO_4[8]\ : OR2
      port map(A => \count_send_time[8]_net_1\, B => N_1145_0, Y
         => count_send_time_e8_0_a2_1_0);
    
    \all_time_write.2.time_already_send[2]\ : DFN1E1C0
      port map(D => un15_time_write, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un7_status_full_ack, Q => 
        \time_already_send[2]\);
    
    \count_send_time[4]\ : DFN1
      port map(D => \count_send_time_RNO[4]_net_1\, CLK => HCLK_c, 
        Q => \count_send_time[4]_net_1\);
    
    \state_RNO[6]\ : OA1C
      port map(A => \send_16_3_time_1_sqmuxa_i_o3_0\, B => N_1027, 
        C => state_tr2_i_0, Y => \state_RNO[6]_net_1\);
    
    \sel_data_0_RNISJ1Q[0]\ : MX2C
      port map(A => N_1327, B => N_1289, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[6]\);
    
    \state_RNIU5T[2]\ : OR2A
      port map(A => N_1030, B => \state[2]_net_1\, Y => 
        time_fifo_ren_1);
    
    \count_send_time[3]\ : DFN1
      port map(D => count_send_time_e3, CLK => HCLK_c, Q => 
        \count_send_time[3]_net_1\);
    
    \count_send_time_RNIKK24_0[20]\ : NOR2
      port map(A => \count_send_time[19]_net_1\, B => 
        \count_send_time[20]_net_1\, Y => state_tr13_0_a2_4);
    
    \sel_data_0_RNIOIAC[0]\ : MX2C
      port map(A => N_1320, B => N_1282, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[13]\);
    
    \count_send_time_RNO_0[29]\ : NOR2A
      port map(A => \count_send_time[28]_net_1\, B => N_1156, Y
         => N_1160);
    
    \count_send_time_RNO[1]\ : OR3C
      port map(A => N_1239, B => N_1237, C => N_1236, Y => 
        count_send_time_e1);
    
    \count_send_time_RNO_1[3]\ : OR3C
      port map(A => \state_0[2]_net_1\, B => 
        \count_send_time[3]_net_1\, C => N_1217, Y => N_1247);
    
    \count_send_time_RNIJPA7[2]\ : NOR2A
      port map(A => \count_send_time[3]_net_1\, B => 
        \count_send_time[2]_net_1\, Y => 
        \state_ns_i_a2_0_a4_0_25_2[5]\);
    
    \count_send_time_RNO_4[20]\ : OR2
      port map(A => \count_send_time[20]_net_1\, B => N_1145_0, Y
         => count_send_time_e20_0_a2_1_0);
    
    \count_send_time_RNO[20]\ : OR3C
      port map(A => N_1107, B => N_1108, C => N_1109, Y => 
        count_send_time_e20);
    
    \state_RNO[7]\ : AO1C
      port map(A => un1_data_send_ok, B => \state[0]_net_1\, C
         => N_1040, Y => \state_RNO[7]_net_1\);
    
    \count_send_time[2]\ : DFN1
      port map(D => count_send_time_e2, CLK => HCLK_c, Q => 
        \count_send_time[2]_net_1\);
    
    \sel_data_RNI955D[0]\ : MX2C
      port map(A => N_1311, B => N_1287, S => \sel_data[0]_net_1\, 
        Y => \data_address[18]\);
    
    \sel_data_0_RNI0MA8_2[0]\ : OR2
      port map(A => \sel_data[1]_net_1\, B => 
        \sel_data_0[0]_net_1\, Y => un27_time_write);
    
    \count_send_time_RNIKK24[20]\ : NOR2B
      port map(A => \count_send_time[19]_net_1\, B => 
        \count_send_time[20]_net_1\, Y => 
        count_send_time_e25_0_o3_m6_0_a2_2);
    
    \state_RNI7PI3[2]\ : OR2B
      port map(A => \state[2]_net_1\, B => HRESETn_c, Y => N_1145);
    
    \count_send_time_RNO_2[10]\ : OR3A
      port map(A => \count_send_time[9]_net_1\, B => N_1225, C
         => count_send_time_e10_0_a2_1_0, Y => N_1273);
    
    \count_send_time_RNO_0[26]\ : OR3A
      port map(A => \count_send_time[25]_net_1\, B => 
        count_send_time_e25_0_o3_N_7_i_0, C => N_1145, Y => 
        N_1163);
    
    \count_send_time_RNO[18]\ : AO1C
      port map(A => \count_send_time[18]_net_1\, B => N_1137, C
         => count_send_time_e18_0_0, Y => count_send_time_e18);
    
    \state_RNO_0[1]\ : NOR3B
      port map(A => \state_0[2]_net_1\, B => state_tr13_0_a2_10, 
        C => state_tr13_0_a2_9, Y => state_tr13_0_a2_14);
    
    \state_RNO_2[1]\ : NOR3A
      port map(A => state_tr13_0_a2_7, B => state_tr13_0_a2_17_0, 
        C => state_tr13_0_a2_17_1, Y => state_tr13_0_a2_12);
    
    \count_send_time_RNI3V2D2[27]\ : OR3B
      port map(A => N_1146, B => \count_send_time[27]_net_1\, C
         => N_1145, Y => N_1156);
    
    \sel_data_0_RNI714P[0]\ : MX2C
      port map(A => N_1279, B => N_1297, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[0]\);
    
    \count_send_time_RNO[6]\ : NOR3A
      port map(A => N_1091, B => N_1253, C => N_1230, Y => 
        \count_send_time_RNO[6]_net_1\);
    
    time_write_RNI6IL9_1 : NOR2A
      port map(A => \time_write\, B => \un20_time_write\, Y => 
        un22_time_write);
    
    \gen_select_address.1.lpp_waveform_dma_selectaddress_I\ : 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I_2\
      port map(nb_burst_available(10) => nb_burst_available(10), 
        nb_burst_available(9) => nb_burst_available(9), 
        nb_burst_available(8) => nb_burst_available(8), 
        nb_burst_available(7) => nb_burst_available(7), 
        nb_burst_available(6) => nb_burst_available(6), 
        nb_burst_available(5) => nb_burst_available(5), 
        nb_burst_available(4) => nb_burst_available(4), 
        nb_burst_available(3) => nb_burst_available(3), 
        nb_burst_available(2) => nb_burst_available(2), 
        nb_burst_available(1) => nb_burst_available(1), 
        nb_burst_available(0) => nb_burst_available(0), 
        status_full_err(1) => status_full_err(1), status_full(1)
         => status_full(1), sel_data(1) => \sel_data[1]_net_1\, 
        sel_data_0(1) => \sel_data_0[1]_net_1\, 
        update_and_sel_5(3) => \update_and_sel_5[3]\, 
        update_and_sel_5(2) => \update_and_sel_5[2]\, 
        addr_data_f1(31) => addr_data_f1(31), addr_data_f1(30)
         => addr_data_f1(30), addr_data_f1(29) => 
        addr_data_f1(29), addr_data_f1(28) => addr_data_f1(28), 
        addr_data_f1(27) => addr_data_f1(27), addr_data_f1(26)
         => addr_data_f1(26), addr_data_f1(25) => 
        addr_data_f1(25), addr_data_f1(24) => addr_data_f1(24), 
        addr_data_f1(23) => addr_data_f1(23), addr_data_f1(22)
         => addr_data_f1(22), addr_data_f1(21) => 
        addr_data_f1(21), addr_data_f1(20) => addr_data_f1(20), 
        addr_data_f1(19) => addr_data_f1(19), addr_data_f1(18)
         => addr_data_f1(18), addr_data_f1(17) => 
        addr_data_f1(17), addr_data_f1(16) => addr_data_f1(16), 
        addr_data_f1(15) => addr_data_f1(15), addr_data_f1(14)
         => addr_data_f1(14), addr_data_f1(13) => 
        addr_data_f1(13), addr_data_f1(12) => addr_data_f1(12), 
        addr_data_f1(11) => addr_data_f1(11), addr_data_f1(10)
         => addr_data_f1(10), addr_data_f1(9) => addr_data_f1(9), 
        addr_data_f1(8) => addr_data_f1(8), addr_data_f1(7) => 
        addr_data_f1(7), addr_data_f1(6) => addr_data_f1(6), 
        addr_data_f1(5) => addr_data_f1(5), addr_data_f1(4) => 
        addr_data_f1(4), addr_data_f1(3) => addr_data_f1(3), 
        addr_data_f1(2) => addr_data_f1(2), addr_data_f1(1) => 
        addr_data_f1(1), addr_data_f1(0) => addr_data_f1(0), 
        status_full_ack(1) => status_full_ack(1), 
        addr_data_vector_94 => \addr_data_vector[126]\, 
        addr_data_vector_91 => \addr_data_vector[123]\, 
        addr_data_vector_89 => \addr_data_vector[121]\, 
        addr_data_vector_87 => \addr_data_vector[119]\, 
        addr_data_vector_86 => \addr_data_vector[118]\, 
        addr_data_vector_85 => \addr_data_vector[117]\, 
        addr_data_vector_84 => \addr_data_vector[116]\, 
        addr_data_vector_83 => \addr_data_vector[115]\, 
        addr_data_vector_67 => \addr_data_vector[99]\, 
        addr_data_vector_66 => \addr_data_vector[98]\, 
        addr_data_vector_65 => \addr_data_vector[97]\, 
        addr_data_vector_64 => \addr_data_vector[96]\, 
        addr_data_vector_75 => \addr_data_vector[107]\, 
        addr_data_vector_73 => \addr_data_vector[105]\, 
        addr_data_vector_81 => \addr_data_vector[113]\, 
        addr_data_vector_79 => \addr_data_vector[111]\, 
        addr_data_vector_77 => \addr_data_vector[109]\, 
        addr_data_vector_24 => \addr_data_vector[56]\, 
        addr_data_vector_31 => \addr_data_vector[63]\, 
        addr_data_vector_16 => \addr_data_vector[48]\, 
        addr_data_vector_14 => \addr_data_vector[46]\, 
        addr_data_vector_18 => \addr_data_vector[50]\, 
        addr_data_vector_26 => \addr_data_vector[58]\, 
        addr_data_vector_29 => \addr_data_vector[61]\, 
        addr_data_vector_28 => \addr_data_vector[60]\, 
        addr_data_vector_5 => \addr_data_vector[37]\, 
        addr_data_vector_4 => \addr_data_vector[36]\, 
        addr_data_vector_6 => \addr_data_vector[38]\, 
        addr_data_vector_12 => \addr_data_vector[44]\, 
        addr_data_vector_10 => \addr_data_vector[42]\, 
        addr_data_vector_7 => \addr_data_vector[39]\, 
        addr_data_vector_8 => \addr_data_vector[40]\, N_913 => 
        N_913, N_910 => N_910, N_908 => N_908, N_906 => N_906, 
        N_905 => N_905, N_904 => N_904, N_903 => N_903, N_902 => 
        N_902, N_1300 => N_1300, N_1299 => N_1299, N_1298 => 
        N_1298, N_1297 => N_1297, N_1294 => N_1294, N_1292 => 
        N_1292, N_1286 => N_1286, N_1284 => N_1284, N_1282 => 
        N_1282, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c);
    
    \count_send_time[24]\ : DFN1
      port map(D => count_send_time_e24, CLK => HCLK_c, Q => 
        \count_send_time[24]_net_1\);
    
    \count_send_time_RNO_1[12]\ : OR2B
      port map(A => \count_send_time[12]_net_1\, B => N_1220, Y
         => N_1080);
    
    \update_RNO[0]\ : OA1
      port map(A => \state[3]_net_1\, B => \state[5]_net_1\, C
         => un1_time_send_ok, Y => update_0_sqmuxa);
    
    \count_send_time_RNO_0[20]\ : AO1B
      port map(A => \count_send_time[19]_net_1\, B => N_1063, C
         => count_send_time_e20_0_a2_0, Y => N_1107);
    
    \sel_data_0_RNICIAC[0]\ : MX2C
      port map(A => N_1317, B => N_1293, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[10]\);
    
    \count_send_time_RNI1RIK1[15]\ : NOR3B
      port map(A => N_1059, B => \count_send_time[15]_net_1\, C
         => N_1145, Y => N_1077);
    
    \count_send_time_RNO[23]\ : OR3C
      port map(A => N_1121, B => N_1122, C => N_1123, Y => 
        count_send_time_e23);
    
    \sel_data_RNI155D[0]\ : MX2C
      port map(A => N_1309, B => N_1285, S => \sel_data[0]_net_1\, 
        Y => \data_address[16]\);
    
    \count_send_time_RNO_1[11]\ : OR2B
      port map(A => \count_send_time[11]_net_1\, B => N_1220, Y
         => N_1169);
    
    \count_send_time_RNO[11]\ : OR3C
      port map(A => N_1167, B => N_1169, C => N_1170, Y => 
        count_send_time_e11);
    
    \count_send_time[27]\ : DFN1
      port map(D => \count_send_time_RNO[27]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[27]_net_1\);
    
    \count_send_time_RNO_1[20]\ : OR2B
      port map(A => \count_send_time[20]_net_1\, B => N_1220, Y
         => N_1108);
    
    \count_send_time_RNO_4[2]\ : AOI1B
      port map(A => \count_send_time[1]_net_1\, B => 
        \count_send_time[0]_net_1\, C => 
        \count_send_time[2]_net_1\, Y => 
        count_send_time_e2_0_a2_0_0);
    
    \count_send_time_RNO_2[20]\ : OR3B
      port map(A => N_1063, B => \count_send_time[19]_net_1\, C
         => count_send_time_e20_0_a2_1_0, Y => N_1109);
    
    \count_send_time_RNO_0[17]\ : OA1C
      port map(A => N_1061, B => N_1145, C => 
        \count_send_time[17]_net_1\, Y => N_1096);
    
    time_select_RNII30M1 : OA1C
      port map(A => N_200, B => N_249, C => \time_select\, Y => 
        \data_ren\);
    
    \sel_data_0_RNIIPAU1[0]\ : OR2A
      port map(A => \data_ren\, B => un27_time_write, Y => 
        data_ren(0));
    
    time_write_RNI6IL9_0 : NOR2A
      port map(A => \time_write\, B => \un13_time_write\, Y => 
        un15_time_write);
    
    \state[3]\ : DFN1C0
      port map(D => \state_RNO_2[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    
    time_fifo_ren : DFN1E0P0
      port map(D => time_fifo_ren_1_i, CLK => HCLK_c, PRE => 
        HRESETn_c, E => \state[0]_net_1\, Q => \time_fifo_ren\);
    
    \count_send_time_RNIK6CT[0]\ : NOR3C
      port map(A => \state_ns_i_a2_0_a4_0_25_1[5]\, B => 
        \state_ns_i_a2_0_a4_0_25_0[5]\, C => 
        \state_ns_i_a2_0_a4_0_25_4[5]\, Y => N_1047_25);
    
    time_write_RNO_0 : OR2
      port map(A => \state[1]_net_1\, B => \state[3]_net_1\, Y
         => un1_state_13_0_a4_0_0);
    
    \count_send_time_RNO_1[1]\ : OR3B
      port map(A => \count_send_time[1]_net_1\, B => 
        \state[2]_net_1\, C => \count_send_time[0]_net_1\, Y => 
        N_1237);
    
    time_select_0 : DFN1E1C0
      port map(D => time_fifo_ren_1, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_816, Q => \time_select_0\);
    
    \sel_data_RNI555D[0]\ : MX2C
      port map(A => N_1310, B => N_1286, S => \sel_data[0]_net_1\, 
        Y => \data_address[17]\);
    
    \count_send_time_RNIJ9211[7]\ : OR3C
      port map(A => N_1223, B => \count_send_time[7]_net_1\, C
         => \count_send_time[8]_net_1\, Y => N_1225);
    
    \count_send_time_RNO_0[18]\ : AOI1B
      port map(A => \count_send_time[18]_net_1\, B => N_1220, C
         => N_1099, Y => count_send_time_e18_0_0);
    
    lpp_dma_send_1word_1 : lpp_dma_send_1word
      port map(Lock => Lock, Request => Request, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, un1_time_send_ok => 
        un1_time_send_ok, time_select => \time_select\, Store => 
        Store, N_1012 => N_1012, Ready => Ready, Fault => Fault, 
        time_send => \time_send\, Grant => Grant);
    
    \all_time_write.0.time_already_send_RNO[0]\ : OR2
      port map(A => status_full_ack(0), B => un29_time_write, Y
         => un17_status_full_ack);
    
    \count_send_time_RNIMBLO1[17]\ : NOR3B
      port map(A => N_1061, B => \count_send_time[17]_net_1\, C
         => N_1145, Y => N_1137);
    
    \count_send_time_RNO_2[31]\ : OR3
      port map(A => N_1161, B => \count_send_time[31]_net_1\, C
         => N_1156, Y => N_1194);
    
    \count_send_time[11]\ : DFN1
      port map(D => count_send_time_e11, CLK => HCLK_c, Q => 
        \count_send_time[11]_net_1\);
    
    \sel_data_RNIQ60E[0]\ : MX2C
      port map(A => N_1315, B => N_905, S => \sel_data[0]_net_1\, 
        Y => \data_address[22]\);
    
    \count_send_time[1]\ : DFN1
      port map(D => count_send_time_e1, CLK => HCLK_c, Q => 
        \count_send_time[1]_net_1\);
    
    \count_send_time[9]\ : DFN1
      port map(D => count_send_time_e9, CLK => HCLK_c, Q => 
        \count_send_time[9]_net_1\);
    
    \sel_data_0_RNI042Q[0]\ : MX2C
      port map(A => N_1328, B => N_1290, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[7]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \count_send_time_RNO_1[8]\ : OR2B
      port map(A => \count_send_time[8]_net_1\, B => N_1220, Y
         => N_1262);
    
    \sel_data_RNIE70E[0]\ : MX2C
      port map(A => N_1306, B => N_910, S => \sel_data[0]_net_1\, 
        Y => \data_address[27]\);
    
    \sel_data_RNIM60E[0]\ : MX2C
      port map(A => N_1314, B => N_904, S => \sel_data[0]_net_1\, 
        Y => \data_address[21]\);
    
    \count_send_time[20]\ : DFN1
      port map(D => count_send_time_e20, CLK => HCLK_c, Q => 
        \count_send_time[20]_net_1\);
    
    \state_ns_i_a2_0_RNO_5[5]\ : NOR2B
      port map(A => state_tr13_0_a2_7, B => state_tr13_0_a2_8, Y
         => \state_ns_i_a2_0_a4_0_19_12[5]\);
    
    \count_send_time[30]\ : DFN1
      port map(D => count_send_time_e30, CLK => HCLK_c, Q => 
        \count_send_time[30]_net_1\);
    
    \count_send_time[15]\ : DFN1
      port map(D => \count_send_time_RNO[15]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[15]_net_1\);
    
    \count_send_time_RNO[16]\ : OA1C
      port map(A => N_1061, B => N_1145_0, C => 
        count_send_time_e16_i_0, Y => 
        \count_send_time_RNO[16]_net_1\);
    
    \DMAWriteFSM_p.sel_data_3_i_a4[1]\ : NOR2A
      port map(A => ready_i_0(3), B => ready_i_0(2), Y => N_1036);
    
    \all_time_write.2.time_already_send_RNISCP08[2]\ : MX2
      port map(A => \time_already_send[3]\, B => 
        \time_already_send[2]\, S => ready_i_0(2), Y => N_1024);
    
    \state_RNO[5]\ : AO1C
      port map(A => N_1026, B => \state[6]_net_1\, C => N_1042, Y
         => \state_RNO[5]_net_1\);
    
    \count_send_time_RNITLAI[4]\ : NOR3B
      port map(A => \count_send_time[3]_net_1\, B => 
        \count_send_time[4]_net_1\, C => N_1217, Y => N_1219);
    
    \count_send_time_RNI7558[13]\ : NOR3A
      port map(A => state_tr13_0_a2_4, B => 
        \count_send_time[18]_net_1\, C => 
        \count_send_time[13]_net_1\, Y => state_tr13_0_a2_9_0);
    
    \count_send_time_RNO_1[18]\ : AO1B
      port map(A => \count_send_time[17]_net_1\, B => N_1061, C
         => count_send_time_e18_0_a2_0_0, Y => N_1099);
    
    \count_send_time_RNIHG24[14]\ : NOR2
      port map(A => \count_send_time[14]_net_1\, B => 
        \count_send_time[15]_net_1\, Y => 
        \state_ns_i_a2_0_a4_0_19_9_0[5]\);
    
    \sel_data_RNI1N0E[0]\ : MX2C
      port map(A => N_1296, B => N_914, S => \sel_data[0]_net_1\, 
        Y => \data_address[31]\);
    
    \count_send_time[18]\ : DFN1
      port map(D => count_send_time_e18, CLK => HCLK_c, Q => 
        \count_send_time[18]_net_1\);
    
    \count_send_time_RNO_0[15]\ : OA1C
      port map(A => N_1059, B => N_1145, C => 
        \count_send_time[15]_net_1\, Y => N_1092);
    
    \count_send_time_RNO[12]\ : OR3C
      port map(A => N_1081, B => N_1080, C => N_1082, Y => 
        count_send_time_e12);
    
    \state[2]\ : DFN1C0
      port map(D => \state_ns_i_a2_0[5]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \state[2]_net_1\);
    
    \count_send_time_RNO_5[30]\ : OR3
      port map(A => N_1075, B => \count_send_time[30]_net_1\, C
         => N_1145_0, Y => count_send_time_e30_0_a2_2_1);
    
    \send_16_3_time[0]\ : DFN1E0P0
      port map(D => \send_16_3_time[2]_net_1\, CLK => HCLK_c, PRE
         => HRESETn_c, E => N_1014, Q => 
        \send_16_3_time[0]_net_1\);
    
    \count_send_time_RNO_3[8]\ : NOR2B
      port map(A => \count_send_time[8]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e8_0_a2_0);
    
    \count_send_time_RNO_0[8]\ : AO1B
      port map(A => \count_send_time[7]_net_1\, B => N_1223, C
         => count_send_time_e8_0_a2_0, Y => N_1260);
    
    \count_send_time_RNO[29]\ : XA1
      port map(A => N_1160, B => \count_send_time[29]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[29]_net_1\);
    
    \count_send_time[6]\ : DFN1
      port map(D => \count_send_time_RNO[6]_net_1\, CLK => HCLK_c, 
        Q => \count_send_time[6]_net_1\);
    
    \send_16_3_time[2]\ : DFN1E0C0
      port map(D => \send_16_3_time[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => N_1014, Q => 
        \send_16_3_time[2]_net_1\);
    
    \state_0[2]\ : DFN1C0
      port map(D => \state_ns_i_a2_0[5]_net_1\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \state_0[2]_net_1\);
    
    \count_send_time_RNIQ858[31]\ : NOR3A
      port map(A => state_tr13_0_a2_2, B => 
        \count_send_time[10]_net_1\, C => 
        \count_send_time[31]_net_1\, Y => state_tr13_0_a2_8);
    
    \count_send_time_RNI089V1[22]\ : OR3B
      port map(A => \count_send_time[21]_net_1\, B => 
        \count_send_time[22]_net_1\, C => N_1066, Y => N_1069);
    
    \state[1]\ : DFN1C0
      port map(D => \state_ns[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[1]_net_1\);
    
    \count_send_time_RNO_4[10]\ : OR2
      port map(A => \count_send_time[10]_net_1\, B => N_1145_0, Y
         => count_send_time_e10_0_a2_1_0);
    
    \count_send_time_RNIRO24[26]\ : OR2
      port map(A => \count_send_time[26]_net_1\, B => 
        \count_send_time[27]_net_1\, Y => state_tr13_0_a2_17_0);
    
    \count_send_time_RNO[17]\ : NOR3A
      port map(A => N_1091, B => N_1096, C => N_1137, Y => 
        \count_send_time_RNO[17]_net_1\);
    
    time_send_RNO_0 : NOR2
      port map(A => \state[2]_net_1\, B => \state[0]_net_1\, Y
         => N_815);
    
    \all_time_write.1.time_already_send_RNI7H7MG[1]\ : MX2
      port map(A => N_1024, B => \time_already_send[1]\, S => 
        ready_i_0(1), Y => N_1025);
    
    \sel_data_RNIT45D[0]\ : MX2C
      port map(A => N_1322, B => N_1284, S => \sel_data[0]_net_1\, 
        Y => \data_address[15]\);
    
    \count_send_time_RNIEPE72[26]\ : NOR3B
      port map(A => \count_send_time[25]_net_1\, B => 
        \count_send_time[26]_net_1\, C => 
        count_send_time_e25_0_o3_N_7_i_0, Y => N_1146);
    
    \state_ns_i_a2_0_RNO_1[5]\ : AOI1B
      port map(A => \state_ns_i_a2_0_a4_0_19_i[5]\, B => 
        \state_0[2]_net_1\, C => N_1050, Y => 
        \state_ns_i_a2_0_0[5]\);
    
    \state_RNO_0[6]\ : OR2B
      port map(A => \send_16_3_time[0]_net_1\, B => 
        \state[7]_net_1\, Y => state_tr2_i_0);
    
    \state_ns_i_a2_0[5]\ : NAND2
      port map(A => N_1049, B => \state_ns_i_a2_0_1[5]\, Y => 
        \state_ns_i_a2_0[5]_net_1\);
    
    \count_send_time_RNO_2[2]\ : OR2B
      port map(A => \count_send_time[2]_net_1\, B => N_1220, Y
         => N_1241);
    
    \count_send_time_RNO_4[24]\ : OR2
      port map(A => \count_send_time[24]_net_1\, B => N_1145_0, Y
         => count_send_time_e24_0_a2_1_0);
    
    \all_time_write.1.time_already_send_RNO[1]\ : OR2
      port map(A => status_full_ack(1), B => un22_time_write, Y
         => un12_status_full_ack);
    
    \state_RNO[3]\ : AO1A
      port map(A => N_1026, B => \state[4]_net_1\, C => N_1033, Y
         => \state_RNO_2[3]\);
    
    \state_RNO[0]\ : AO1
      port map(A => \state[0]_net_1\, B => un1_data_send_ok, C
         => \state[1]_net_1\, Y => \state_RNO_1[0]\);
    
    \state_ns_i_a2_0_RNO[5]\ : AND2
      port map(A => N_1048, B => \state_ns_i_a2_0_0[5]\, Y => 
        \state_ns_i_a2_0_1[5]\);
    
    \sel_data_0_RNIKJ0Q[0]\ : MX2C
      port map(A => N_1325, B => N_1301, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[4]\);
    
    \count_send_time_RNO_2[13]\ : OR3
      port map(A => N_1145, B => \count_send_time[13]_net_1\, C
         => N_1057, Y => N_1087);
    
    \state_RNO_1[1]\ : NOR3C
      port map(A => state_tr13_0_a2_9_0, B => state_tr13_0_a2_8, 
        C => state_tr13_0_a2_12, Y => state_tr13_0_a2_15);
    
    \state_ns_i_a2_0_RNO_4[5]\ : OR2B
      port map(A => \state[3]_net_1\, B => un1_time_send_ok, Y
         => N_1050);
    
    \count_send_time_RNO_0[4]\ : OR3A
      port map(A => \count_send_time[3]_net_1\, B => N_1217, C
         => N_1145, Y => N_1227);
    
    \count_send_time_RNIL0C32[15]\ : OR3C
      port map(A => N_1059, B => \count_send_time[15]_net_1\, C
         => count_send_time_e25_0_o3_m6_0_a2_7, Y => 
        count_send_time_e25_0_o3_N_7_i_0);
    
    \sel_data_RNI270E[0]\ : MX2C
      port map(A => N_1303, B => N_907, S => \sel_data[0]_net_1\, 
        Y => \data_address[24]\);
    
    \count_send_time_RNO_1[31]\ : OR2B
      port map(A => \count_send_time[31]_net_1\, B => N_1220, Y
         => N_1193);
    
    time_fifo_ren_RNIGHOH : OR2A
      port map(A => \time_ren\, B => \un20_time_write\, Y => 
        time_ren(1));
    
    \count_send_time_RNO_0[5]\ : OR2A
      port map(A => N_1219, B => N_1145, Y => N_1228);
    
    \count_send_time_RNO_3[30]\ : NOR2B
      port map(A => \count_send_time[30]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e30_0_a2_0_0);
    
    \count_send_time_RNO_0[23]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[23]_net_1\, C => N_1069, Y => N_1121);
    
    \count_send_time_RNO_0[24]\ : AO1C
      port map(A => N_1069, B => \count_send_time[23]_net_1\, C
         => count_send_time_e24_0_a2_0_0, Y => N_1173);
    
    time_send : DFN1E1C0
      port map(D => time_send_0_sqmuxa, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_815, Q => \time_send\);
    
    \count_send_time_RNO_0[31]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[31]_net_1\, C => N_1162, Y => N_1191);
    
    time_select_RNIIPAU1 : OR2A
      port map(A => \data_ren\, B => \un13_time_write\, Y => 
        data_ren(2));
    
    \count_send_time_RNO_3[10]\ : NOR2B
      port map(A => \count_send_time[10]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e10_0_a2_0);
    
    \count_send_time_RNO_0[1]\ : OR3A
      port map(A => \count_send_time[0]_net_1\, B => 
        \count_send_time[1]_net_1\, C => N_1145_0, Y => N_1239);
    
    \update[0]\ : DFN1E0C0
      port map(D => update_0_sqmuxa, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un1_state_12, Q => \update[0]_net_1\);
    
    \count_send_time_RNO_1[23]\ : OR2B
      port map(A => \count_send_time[23]_net_1\, B => N_1220, Y
         => N_1122);
    
    \count_send_time_RNO[28]\ : XA1A
      port map(A => N_1156, B => \count_send_time[28]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[28]_net_1\);
    
    \count_send_time_RNO_2[23]\ : OR3
      port map(A => N_1145_0, B => \count_send_time[23]_net_1\, C
         => N_1069, Y => N_1123);
    
    \count_send_time_RNO_1[24]\ : OR2B
      port map(A => \count_send_time[24]_net_1\, B => N_1220, Y
         => N_1172);
    
    \count_send_time_RNIBG24[12]\ : NOR2
      port map(A => \count_send_time[11]_net_1\, B => 
        \count_send_time[12]_net_1\, Y => state_tr13_0_a2_2);
    
    \count_send_time_RNO_2[24]\ : OR3A
      port map(A => \count_send_time[23]_net_1\, B => N_1069, C
         => count_send_time_e24_0_a2_1_0, Y => N_1175);
    
    \count_send_time[23]\ : DFN1
      port map(D => count_send_time_e23, CLK => HCLK_c, Q => 
        \count_send_time[23]_net_1\);
    
    \count_send_time[22]\ : DFN1
      port map(D => count_send_time_e22, CLK => HCLK_c, Q => 
        \count_send_time[22]_net_1\);
    
    \state_ns_i_a2_0_RNO_6[5]\ : NOR3
      port map(A => state_tr13_0_a2_17_0, B => 
        state_tr13_0_a2_17_1, C => state_tr13_0_a2_9, Y => 
        \state_ns_i_a2_0_a4_0_19_11[5]\);
    
    \sel_data_RNII60E[0]\ : MX2C
      port map(A => N_1313, B => N_903, S => \sel_data[0]_net_1\, 
        Y => \data_address[20]\);
    
    \update_RNIOECD_2[0]\ : OR2A
      port map(A => \update[0]_net_1\, B => un27_time_write, Y
         => \update_and_sel_7[0]\);
    
    \count_send_time_RNO_4[22]\ : OR2
      port map(A => \count_send_time[22]_net_1\, B => N_1145_0, Y
         => count_send_time_e22_0_a2_1_0);
    
    \count_send_time[16]\ : DFN1
      port map(D => \count_send_time_RNO[16]_net_1\, CLK => 
        HCLK_c, Q => \count_send_time[16]_net_1\);
    
    \count_send_time_RNIHPUE1[14]\ : NOR3B
      port map(A => \count_send_time[13]_net_1\, B => 
        \count_send_time[14]_net_1\, C => N_1057, Y => N_1059);
    
    \count_send_time_RNO[30]\ : OR3C
      port map(A => N_1126, B => count_send_time_e30_0_0, C => 
        N_1128, Y => count_send_time_e30);
    
    \count_send_time_RNO[21]\ : OR3C
      port map(A => N_1112, B => N_1113, C => N_1114, Y => 
        count_send_time_e21);
    
    \sel_data_0_RNIGHOH[0]\ : OR2A
      port map(A => \time_ren\, B => un27_time_write, Y => 
        time_ren(0));
    
    \count_send_time_RNO_2[12]\ : OR3A
      port map(A => \count_send_time[11]_net_1\, B => N_1159, C
         => count_send_time_e12_0_a2_1_0, Y => N_1082);
    
    \all_time_write.2.time_already_send_RNO[2]\ : OR2
      port map(A => status_full_ack(2), B => un15_time_write, Y
         => un7_status_full_ack);
    
    \all_time_write.1.time_already_send[1]\ : DFN1E1C0
      port map(D => un22_time_write, CLK => HCLK_c, CLR => 
        HRESETn_c, E => un12_status_full_ack, Q => 
        \time_already_send[1]\);
    
    \gen_select_address.3.lpp_waveform_dma_selectaddress_I\ : 
        \lpp_waveform_dma_selectaddress_gen_select_address.3.lpp_waveform_dma_selectaddress_I\
      port map(nb_burst_available(10) => nb_burst_available(10), 
        nb_burst_available(9) => nb_burst_available(9), 
        nb_burst_available(8) => nb_burst_available(8), 
        nb_burst_available(7) => nb_burst_available(7), 
        nb_burst_available(6) => nb_burst_available(6), 
        nb_burst_available(5) => nb_burst_available(5), 
        nb_burst_available(4) => nb_burst_available(4), 
        nb_burst_available(3) => nb_burst_available(3), 
        nb_burst_available(2) => nb_burst_available(2), 
        nb_burst_available(1) => nb_burst_available(1), 
        nb_burst_available(0) => nb_burst_available(0), 
        status_full_err(3) => status_full_err(3), status_full(3)
         => status_full(3), sel_data(1) => \sel_data[1]_net_1\, 
        sel_data_0(1) => \sel_data_0[1]_net_1\, 
        update_and_sel_1(7) => \update_and_sel_1[7]\, 
        update_and_sel_1(6) => \update_and_sel_1[6]\, 
        addr_data_f3(31) => addr_data_f3(31), addr_data_f3(30)
         => addr_data_f3(30), addr_data_f3(29) => 
        addr_data_f3(29), addr_data_f3(28) => addr_data_f3(28), 
        addr_data_f3(27) => addr_data_f3(27), addr_data_f3(26)
         => addr_data_f3(26), addr_data_f3(25) => 
        addr_data_f3(25), addr_data_f3(24) => addr_data_f3(24), 
        addr_data_f3(23) => addr_data_f3(23), addr_data_f3(22)
         => addr_data_f3(22), addr_data_f3(21) => 
        addr_data_f3(21), addr_data_f3(20) => addr_data_f3(20), 
        addr_data_f3(19) => addr_data_f3(19), addr_data_f3(18)
         => addr_data_f3(18), addr_data_f3(17) => 
        addr_data_f3(17), addr_data_f3(16) => addr_data_f3(16), 
        addr_data_f3(15) => addr_data_f3(15), addr_data_f3(14)
         => addr_data_f3(14), addr_data_f3(13) => 
        addr_data_f3(13), addr_data_f3(12) => addr_data_f3(12), 
        addr_data_f3(11) => addr_data_f3(11), addr_data_f3(10)
         => addr_data_f3(10), addr_data_f3(9) => addr_data_f3(9), 
        addr_data_f3(8) => addr_data_f3(8), addr_data_f3(7) => 
        addr_data_f3(7), addr_data_f3(6) => addr_data_f3(6), 
        addr_data_f3(5) => addr_data_f3(5), addr_data_f3(4) => 
        addr_data_f3(4), addr_data_f3(3) => addr_data_f3(3), 
        addr_data_f3(2) => addr_data_f3(2), addr_data_f3(1) => 
        addr_data_f3(1), addr_data_f3(0) => addr_data_f3(0), 
        status_full_ack(3) => status_full_ack(3), 
        addr_data_vector_61 => \addr_data_vector[97]\, 
        addr_data_vector_60 => \addr_data_vector[96]\, 
        addr_data_vector_27 => \addr_data_vector[63]\, 
        addr_data_vector_25 => \addr_data_vector[61]\, 
        addr_data_vector_24 => \addr_data_vector[60]\, 
        addr_data_vector_22 => \addr_data_vector[58]\, 
        addr_data_vector_20 => \addr_data_vector[56]\, 
        addr_data_vector_0 => \addr_data_vector[36]\, 
        addr_data_vector_6 => \addr_data_vector[42]\, 
        addr_data_vector_4 => \addr_data_vector[40]\, 
        addr_data_vector_3 => \addr_data_vector[39]\, 
        addr_data_vector_2 => \addr_data_vector[38]\, 
        addr_data_vector_1 => \addr_data_vector[37]\, 
        addr_data_vector_14 => \addr_data_vector[50]\, 
        addr_data_vector_12 => \addr_data_vector[48]\, 
        addr_data_vector_10 => \addr_data_vector[46]\, 
        addr_data_vector_8 => \addr_data_vector[44]\, 
        addr_data_vector_63 => \addr_data_vector[99]\, 
        addr_data_vector_90 => \addr_data_vector[126]\, 
        addr_data_vector_87 => \addr_data_vector[123]\, 
        addr_data_vector_85 => \addr_data_vector[121]\, 
        addr_data_vector_62 => \addr_data_vector[98]\, 
        addr_data_vector_69 => \addr_data_vector[105]\, 
        addr_data_vector_73 => \addr_data_vector[109]\, 
        addr_data_vector_71 => \addr_data_vector[107]\, 
        addr_data_vector_77 => \addr_data_vector[113]\, 
        addr_data_vector_79 => \addr_data_vector[115]\, 
        addr_data_vector_82 => \addr_data_vector[118]\, 
        addr_data_vector_83 => \addr_data_vector[119]\, 
        addr_data_vector_75 => \addr_data_vector[111]\, 
        addr_data_vector_80 => \addr_data_vector[116]\, 
        addr_data_vector_81 => \addr_data_vector[117]\, N_914 => 
        N_914, N_912 => N_912, N_911 => N_911, N_909 => N_909, 
        N_907 => N_907, N_1301 => N_1301, N_1293 => N_1293, 
        N_1291 => N_1291, N_1290 => N_1290, N_1289 => N_1289, 
        N_1288 => N_1288, N_1287 => N_1287, N_1285 => N_1285, 
        N_1283 => N_1283, N_1281 => N_1281, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    \state_ns_i_a2_0_RNO_7[5]\ : NOR3C
      port map(A => state_tr13_0_a2_10, B => state_tr13_0_a2_9_0, 
        C => N_1047_25, Y => \state_ns_i_a2_0_a4_0_19_15[5]\);
    
    \count_send_time_RNO_2[11]\ : OR3
      port map(A => N_1145_0, B => \count_send_time[11]_net_1\, C
         => N_1159, Y => N_1170);
    
    \count_send_time_RNO[5]\ : XA1A
      port map(A => N_1228, B => \count_send_time[5]_net_1\, C
         => N_1091, Y => \count_send_time_RNO[5]_net_1\);
    
    \count_send_time[19]\ : DFN1
      port map(D => count_send_time_e19, CLK => HCLK_c, Q => 
        \count_send_time[19]_net_1\);
    
    \count_send_time_RNO_3[20]\ : NOR2B
      port map(A => \count_send_time[20]_net_1\, B => 
        \state_0[2]_net_1\, Y => count_send_time_e20_0_a2_0);
    
    \sel_data_0_RNICI8P[0]\ : MX2C
      port map(A => N_1316, B => N_1292, S => 
        \sel_data_0[0]_net_1\, Y => \data_address[9]\);
    
    \count_send_time_RNO_0[22]\ : AO1C
      port map(A => N_1066, B => \count_send_time[21]_net_1\, C
         => count_send_time_e22_0_a2_0, Y => N_1117);
    
    \count_send_time_RNO[15]\ : NOR3A
      port map(A => N_1091, B => N_1092, C => N_1077, Y => 
        \count_send_time_RNO[15]_net_1\);
    
    \count_send_time_RNO_0[21]\ : OR3C
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[21]_net_1\, C => N_1066, Y => N_1112);
    
    \count_send_time_RNO_1[22]\ : OR2B
      port map(A => \count_send_time[22]_net_1\, B => N_1220, Y
         => N_1118);
    
    \update_RNIPECD_1[1]\ : NOR2A
      port map(A => \update[1]_net_1\, B => \un13_time_write\, Y
         => \update_and_sel_3[5]\);
    
    \count_send_time_RNO_2[22]\ : OR3A
      port map(A => \count_send_time[21]_net_1\, B => N_1066, C
         => count_send_time_e22_0_a2_1_0, Y => N_1119);
    
    \state_0_RNIAU89[2]\ : OR2B
      port map(A => \state_0[2]_net_1\, B => HRESETn_c, Y => 
        N_1145_0);
    
    \state_RNI8UM1[0]\ : AO1B
      port map(A => \state[0]_net_1\, B => un1_data_send_ok, C
         => N_1030, Y => un1_state_12);
    
    DMA2AHB_1 : DMA2AHB
      port map(hburst_c(2) => hburst_c(2), hburst_c(1) => 
        hburst_c(1), hburst_c(0) => hburst_c(0), htrans_c(1) => 
        htrans_c(1), htrans_c(0) => htrans_c(0), un7_dmain(66)
         => \un7_dmain[66]\, hsize_c(1) => hsize_c(1), hsize_c(0)
         => hsize_c(0), AHB_Master_In_c_5 => AHB_Master_In_c_5, 
        AHB_Master_In_c_4 => AHB_Master_In_c_4, AHB_Master_In_c_0
         => AHB_Master_In_c_0, AHB_Master_In_c_3 => 
        AHB_Master_In_c_3, haddr_c(31) => haddr_c(31), 
        haddr_c(30) => haddr_c(30), haddr_c(29) => haddr_c(29), 
        haddr_c(28) => haddr_c(28), haddr_c(27) => haddr_c(27), 
        haddr_c(26) => haddr_c(26), haddr_c(25) => haddr_c(25), 
        haddr_c(24) => haddr_c(24), haddr_c(23) => haddr_c(23), 
        haddr_c(22) => haddr_c(22), haddr_c(21) => haddr_c(21), 
        haddr_c(20) => haddr_c(20), haddr_c(19) => haddr_c(19), 
        haddr_c(18) => haddr_c(18), haddr_c(17) => haddr_c(17), 
        haddr_c(16) => haddr_c(16), haddr_c(15) => haddr_c(15), 
        haddr_c(14) => haddr_c(14), haddr_c(13) => haddr_c(13), 
        haddr_c(12) => haddr_c(12), haddr_c(11) => haddr_c(11), 
        haddr_c(10) => haddr_c(10), haddr_c(9) => haddr_c(9), 
        haddr_c(8) => haddr_c(8), haddr_c(7) => haddr_c(7), 
        haddr_c(6) => haddr_c(6), haddr_c(5) => haddr_c(5), 
        haddr_c(4) => haddr_c(4), haddr_c(3) => haddr_c(3), 
        haddr_c(2) => haddr_c(2), haddr_c(1) => haddr_c(1), 
        haddr_c(0) => haddr_c(0), hwrite_c => hwrite_c, Ready => 
        Ready, N_1012 => N_1012, Grant => Grant, 
        IdlePhase_RNI03G71 => IdlePhase_RNI03G71, OKAY => OKAY, 
        Fault => Fault, N_1011 => N_1011, N_1013 => N_1013, N_43
         => N_43, time_select_0 => \time_select_0\, N_960 => 
        N_960, N_959 => N_959, N_958 => N_958, N_957 => N_957, 
        N_964 => N_964, N_963 => N_963, N_962 => N_962, N_961 => 
        N_961, N_955 => N_955, N_954 => N_954, N_953 => N_953, 
        N_952 => N_952, N_951 => N_951, N_950 => N_950, N_949 => 
        N_949, N_948 => N_948, N_947 => N_947, N_956 => N_956, 
        N_965 => N_965, N_966 => N_966, N_967 => N_967, N_968 => 
        N_968, N_969 => N_969, N_970 => N_970, N_971 => N_971, 
        N_972 => N_972, N_973 => N_973, N_974 => N_974, N_975 => 
        N_975, N_976 => N_976, N_977 => N_977, HRESETn_c => 
        HRESETn_c, N_978 => N_978, HCLK_c => HCLK_c);
    
    \count_send_time_RNO_1[21]\ : OR2B
      port map(A => \count_send_time[21]_net_1\, B => N_1220, Y
         => N_1113);
    
    \count_send_time_RNO_0[19]\ : OR3B
      port map(A => \state[2]_net_1\, B => 
        \count_send_time[19]_net_1\, C => N_1063, Y => N_1103);
    
    \count_send_time_RNIVO24[29]\ : OR2B
      port map(A => \count_send_time[29]_net_1\, B => 
        \count_send_time[28]_net_1\, Y => N_1075);
    
    \count_send_time_RNO_2[21]\ : OR3
      port map(A => N_1145, B => \count_send_time[21]_net_1\, C
         => N_1066, Y => N_1114);
    
    \count_send_time_RNO[9]\ : OR3C
      port map(A => N_1265, B => N_1267, C => N_1268, Y => 
        count_send_time_e9);
    
    \state_ns_i_a2_0_RNO_0[5]\ : AO1C
      port map(A => N_1027, B => \send_16_3_time_1_sqmuxa_i_o3_0\, 
        C => \state_ns_i_a2_0_a3_0[5]_net_1\, Y => N_1048);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform_fifo_arbiter is

    port( wdata       : out   std_logic_vector(31 downto 0);
          data_wen    : out   std_logic_vector(3 downto 0);
          valid_ack   : out   std_logic_vector(3 downto 0);
          time_wen    : out   std_logic_vector(3 downto 0);
          data_f3_out : in    std_logic_vector(159 downto 64);
          data_f2_out : in    std_logic_vector(159 downto 64);
          data_f1_out : in    std_logic_vector(159 downto 64);
          data_f0_out : in    std_logic_vector(159 downto 64);
          valid_out_i : in    std_logic_vector(1 to 1);
          ready_i_0   : in    std_logic_vector(3 downto 0);
          valid_out_3 : in    std_logic;
          valid_out_2 : in    std_logic;
          valid_out_0 : in    std_logic;
          HRESETn_c   : in    std_logic;
          HCLK_c      : in    std_logic
        );

end lpp_waveform_fifo_arbiter;

architecture DEF_ARCH of lpp_waveform_fifo_arbiter is 

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \data_valid_and_ready_3[0]_net_1\, 
        \data_valid_and_ready_2[0]_net_1\, 
        \data_valid_and_ready_1[0]_net_1\, 
        \data_valid_and_ready_0[0]_net_1\, 
        \data_valid_and_ready_3[2]_net_1\, 
        \data_valid_and_ready_2[2]_net_1\, 
        \data_valid_and_ready_1[2]_net_1\, 
        \data_valid_and_ready_0[2]_net_1\, N_863_2, 
        \state[4]_net_1\, \data_temp_5_i_a2_0_0[32]_net_1\, 
        N_1580_0, N_863_1, N_863_0, N_1580_3, 
        \data_valid_and_ready[1]_net_1\, N_1580_2, N_1580_1, 
        \state_0[4]\, N_860_i, N_860, \time_wen_3_i[0]\, 
        \time_wen_3[0]\, N_859_i, N_859, N_857_i, N_857, 
        state_0_sqmuxa_i_i, state_0_sqmuxa_i, 
        \data_temp_5_i_0[32]\, N_912_i, N_769, N_864, 
        \data_temp_5_i_0[33]\, N_770, N_867, 
        \data_temp_5_i_0[34]\, N_848, N_870, 
        \data_temp_5_i_0[35]\, N_849, N_873, 
        \data_temp_5_i_0[36]\, N_850, N_1650, 
        \data_temp_5_i_0[37]\, N_851, N_1653, 
        \data_temp_5_i_0[38]\, N_852, N_1656, 
        \data_temp_5_i_0[39]\, N_853, N_1659, 
        \data_temp_5_i_0[40]\, N_854, N_1662, 
        \data_temp_5_i_0[41]\, N_841, N_1665, 
        \data_temp_5_i_0[42]\, N_842, N_1668, 
        \data_temp_5_i_0[43]\, N_843, N_897, 
        \data_temp_5_i_0[92]\, N_794, N_900, 
        \data_temp_5_i_0[93]\, N_795, N_902, 
        \data_temp_5_i_0[124]\, N_1681, N_904, 
        \data_temp_5_i_0[125]\, N_1682, N_906, 
        \data_temp_5_i_0[91]\, N_793, N_908, 
        \data_temp_5_i_0[123]\, N_1680, N_910, 
        \time_wen_3_i_a2_0[3]_net_1\, 
        \data_valid_and_ready[3]_net_1\, \state_ns_i_i_a2_1[0]\, 
        \state[2]_net_1\, \state[1]_net_1\, \state[3]_net_1\, 
        N_239, N_898, N_237, N_1669, N_235, N_1666, N_233, N_1663, 
        N_231, N_1660, N_229, N_1657, N_227, N_1654, N_225, 
        N_1651, N_223, N_874, N_221, N_871, N_219, N_868, N_215, 
        N_865, N_251, N_913, N_249, N_247, N_914, N_245, N_915, 
        N_243, N_241, N_863, N_861, N_1306, \state[0]_net_1\, 
        N_917, N_858, \data_temp[64]_net_1\, N_1685, 
        \data_temp[65]_net_1\, N_1686, \data_temp[66]_net_1\, 
        N_1687, \data_temp[67]_net_1\, N_1688, 
        \data_temp[68]_net_1\, N_1689, \data_temp[69]_net_1\, 
        N_762, \data_temp[70]_net_1\, N_763, 
        \data_temp[71]_net_1\, N_764, \data_temp[72]_net_1\, 
        N_765, \data_temp[73]_net_1\, N_766, 
        \data_temp[74]_net_1\, N_767, \data_temp[75]_net_1\, 
        N_768, N_1731, N_1718, N_1693, N_1694, N_1730, N_1692, 
        \data_temp[123]_net_1\, \data_temp[125]_net_1\, 
        \data_temp[124]_net_1\, N_916, N_1580, N_1675, N_1676, 
        N_1677, N_1678, N_1679, N_1683, N_1684, N_1690, N_1691, 
        N_1695, N_1696, N_1697, N_1698, N_1699, N_1700, N_1701, 
        N_1702, N_1703, N_1704, N_1705, N_1706, N_1707, N_1708, 
        N_1709, N_1710, N_1711, N_1712, N_1713, N_1714, N_1715, 
        N_1716, N_1717, N_1719, N_1720, N_1721, N_1722, N_1723, 
        N_1724, N_1725, N_1726, N_1727, N_1728, N_1729, N_1732, 
        N_1733, N_1734, N_1735, N_1736, N_1737, N_1738, N_1739, 
        N_1740, N_729, N_730, N_731, N_732, N_733, N_734, N_735, 
        N_736, N_737, N_738, N_739, N_740, N_741, N_742, N_743, 
        N_744, N_745, N_746, N_747, N_748, N_749, N_750, N_751, 
        N_752, \data_valid_and_ready[2]_net_1\, N_753, N_754, 
        N_755, N_756, N_757, N_758, N_759, N_760, N_761, N_771, 
        N_772, N_773, N_774, N_775, N_776, N_777, N_778, N_779, 
        N_780, N_781, N_782, N_783, N_784, N_785, N_786, N_787, 
        N_788, N_789, N_790, N_791, N_792, N_796, N_797, N_798, 
        N_799, N_800, N_801, N_802, N_803, N_804, N_805, N_806, 
        N_807, N_808, N_809, N_810, N_811, N_812, N_813, N_814, 
        N_815, N_816, N_817, N_818, N_819, N_820, N_821, N_822, 
        N_823, N_824, N_825, N_826, N_827, N_828, N_829, N_830, 
        N_831, N_832, N_833, N_834, N_835, N_836, 
        \data_valid_and_ready[0]_net_1\, N_837, N_838, N_839, 
        N_840, N_844, N_845, N_846, N_847, \data_wen_3[0]\, 
        \time_en_temp[0]_net_1\, \data_wen_3[2]\, 
        \time_en_temp[2]_net_1\, \data_wen_3[3]\, 
        \time_en_temp[3]_net_1\, \data_selected[127]\, 
        \data_selected[159]\, N_696, \data_temp[127]_net_1\, 
        N_728, \data_temp_5[95]\, \data_temp_5[127]\, 
        \data_temp_5[14]\, \data_temp[46]_net_1\, 
        \data_temp_5[13]\, \data_temp[45]_net_1\, 
        \data_temp_5[12]\, \data_temp[44]_net_1\, 
        \data_temp_5[11]\, \data_temp[43]_net_1\, 
        \data_temp_5[10]\, \data_temp[42]_net_1\, 
        \data_temp_5[9]\, \data_temp[41]_net_1\, \data_temp_5[8]\, 
        \data_temp[40]_net_1\, \data_temp_5[7]\, 
        \data_temp[39]_net_1\, \data_temp_5[6]\, 
        \data_temp[38]_net_1\, \data_temp_5[5]\, 
        \data_temp[37]_net_1\, \data_temp_5[4]\, 
        \data_temp[36]_net_1\, \data_temp_5[3]\, 
        \data_temp[35]_net_1\, \data_temp_5[2]\, 
        \data_temp[34]_net_1\, \data_temp_5[1]\, 
        \data_temp[33]_net_1\, \data_temp_5[0]\, 
        \data_temp[32]_net_1\, \data_5[31]\, 
        \data_temp[31]_net_1\, \data_5[30]\, 
        \data_temp[30]_net_1\, \data_5[29]\, 
        \data_temp[29]_net_1\, \data_5[28]\, 
        \data_temp[28]_net_1\, \data_5[27]\, 
        \data_temp[27]_net_1\, \data_5[26]\, 
        \data_temp[26]_net_1\, \data_5[25]\, 
        \data_temp[25]_net_1\, \data_5[24]\, 
        \data_temp[24]_net_1\, \data_5[23]\, 
        \data_temp[23]_net_1\, \data_5[22]\, 
        \data_temp[22]_net_1\, \data_5[21]\, 
        \data_temp[21]_net_1\, \data_5[20]\, 
        \data_temp[20]_net_1\, \data_5[19]\, 
        \data_temp[19]_net_1\, \data_5[18]\, 
        \data_temp[18]_net_1\, \data_5[17]\, 
        \data_temp[17]_net_1\, \data_5[16]\, 
        \data_temp[16]_net_1\, \data_5[15]\, 
        \data_temp[15]_net_1\, \data_5[14]\, 
        \data_temp[14]_net_1\, \data_5[13]\, 
        \data_temp[13]_net_1\, \data_5[12]\, 
        \data_temp[12]_net_1\, \data_5[11]\, 
        \data_temp[11]_net_1\, \data_5[10]\, 
        \data_temp[10]_net_1\, \data_5[9]\, \data_temp[9]_net_1\, 
        \data_5[8]\, \data_temp[8]_net_1\, \data_5[7]\, 
        \data_temp[7]_net_1\, \data_5[6]\, \data_temp[6]_net_1\, 
        \data_selected[76]\, \data_selected[77]\, 
        \data_selected[78]\, \data_selected[79]\, 
        \data_selected[126]\, \data_selected[158]\, N_645, 
        \data_temp[76]_net_1\, N_646, \data_temp[77]_net_1\, 
        N_647, \data_temp[78]_net_1\, N_648, 
        \data_temp[79]_net_1\, N_695, \data_temp[126]_net_1\, 
        N_727, \data_temp_5[44]\, \data_temp_5[45]\, 
        \data_temp_5[46]\, \data_temp_5[47]\, \data_temp_5[94]\, 
        \data_temp_5[126]\, \data_temp_5[31]\, 
        \data_temp[63]_net_1\, \data_temp_5[30]\, 
        \data_temp[62]_net_1\, \data_temp_5[29]\, 
        \data_temp[61]_net_1\, \data_temp_5[28]\, 
        \data_temp[60]_net_1\, \data_temp_5[27]\, 
        \data_temp[59]_net_1\, \data_temp_5[26]\, 
        \data_temp[58]_net_1\, \data_temp_5[25]\, 
        \data_temp[57]_net_1\, \data_temp_5[24]\, 
        \data_temp[56]_net_1\, \data_temp_5[23]\, 
        \data_temp[55]_net_1\, \data_temp_5[22]\, 
        \data_temp[54]_net_1\, \data_temp_5[21]\, 
        \data_temp[53]_net_1\, \data_temp_5[20]\, 
        \data_temp[52]_net_1\, \data_temp_5[19]\, 
        \data_temp[51]_net_1\, \data_temp_5[18]\, 
        \data_temp[50]_net_1\, \data_temp_5[17]\, 
        \data_temp[49]_net_1\, \data_temp_5[16]\, 
        \data_temp[48]_net_1\, \data_temp_5[15]\, 
        \data_temp[47]_net_1\, N_928, N_929, \data_selected[80]\, 
        \data_selected[81]\, \data_selected[82]\, 
        \data_selected[83]\, \data_selected[84]\, 
        \data_selected[85]\, \data_selected[86]\, 
        \data_selected[87]\, \data_selected[88]\, 
        \data_selected[89]\, \data_selected[90]\, 
        \data_selected[91]\, \data_selected[92]\, 
        \data_selected[93]\, \data_selected[94]\, 
        \data_selected[95]\, \data_selected[112]\, 
        \data_selected[144]\, N_649, \data_temp[80]_net_1\, N_650, 
        \data_temp[81]_net_1\, N_651, \data_temp[82]_net_1\, 
        N_652, \data_temp[83]_net_1\, N_653, 
        \data_temp[84]_net_1\, N_654, \data_temp[85]_net_1\, 
        N_655, \data_temp[86]_net_1\, N_656, 
        \data_temp[87]_net_1\, N_657, \data_temp[88]_net_1\, 
        N_658, \data_temp[89]_net_1\, N_659, 
        \data_temp[90]_net_1\, N_660, \data_temp[91]_net_1\, 
        N_661, \data_temp[92]_net_1\, N_662, 
        \data_temp[93]_net_1\, N_663, \data_temp[94]_net_1\, 
        N_664, \data_temp[95]_net_1\, N_681, 
        \data_temp[112]_net_1\, N_713, \data_temp_5[48]\, 
        \data_temp_5[49]\, \data_temp_5[50]\, \data_temp_5[51]\, 
        \data_temp_5[52]\, \data_temp_5[53]\, \data_temp_5[54]\, 
        \data_temp_5[55]\, \data_temp_5[56]\, \data_temp_5[57]\, 
        \data_temp_5[58]\, \data_temp_5[59]\, \data_temp_5[60]\, 
        \data_temp_5[61]\, \data_temp_5[62]\, \data_temp_5[63]\, 
        \data_temp_5[80]\, \data_temp_5[112]\, \data_5[5]\, 
        \data_temp[5]_net_1\, \data_5[4]\, \data_temp[4]_net_1\, 
        \data_5[3]\, \data_temp[3]_net_1\, \data_5[2]\, 
        \data_temp[2]_net_1\, \data_5[1]\, \data_temp[1]_net_1\, 
        \data_5[0]\, \data_temp[0]_net_1\, \data_selected[108]\, 
        \data_selected[110]\, \data_selected[140]\, 
        \data_selected[142]\, N_677, \data_temp[108]_net_1\, 
        N_679, \data_temp[110]_net_1\, N_709, N_711, 
        \data_temp_5[76]\, \data_temp_5[78]\, \data_temp_5[108]\, 
        \data_temp_5[110]\, \data_selected[107]\, 
        \data_selected[111]\, \data_selected[139]\, 
        \data_selected[143]\, N_676, \data_temp[107]_net_1\, 
        N_680, \data_temp[111]_net_1\, N_708, N_712, 
        \data_temp_5[75]\, \data_temp_5[79]\, \data_temp_5[107]\, 
        \data_temp_5[111]\, \data_selected[106]\, 
        \data_selected[113]\, \data_selected[138]\, 
        \data_selected[145]\, N_675, \data_temp[106]_net_1\, 
        N_682, \data_temp[113]_net_1\, N_707, N_714, 
        \data_temp_5[74]\, \data_temp_5[81]\, \data_temp_5[106]\, 
        \data_temp_5[113]\, \data_selected[105]\, 
        \data_selected[114]\, \data_selected[137]\, 
        \data_selected[146]\, N_674, \data_temp[105]_net_1\, 
        N_683, \data_temp[114]_net_1\, N_706, N_715, 
        \data_temp_5[73]\, \data_temp_5[82]\, \data_temp_5[105]\, 
        \data_temp_5[114]\, \data_selected[104]\, 
        \data_selected[115]\, \data_selected[136]\, 
        \data_selected[147]\, N_673, \data_temp[104]_net_1\, 
        N_684, \data_temp[115]_net_1\, N_705, N_716, 
        \data_temp_5[72]\, \data_temp_5[83]\, \data_temp_5[104]\, 
        \data_temp_5[115]\, \data_selected[103]\, 
        \data_selected[116]\, \data_selected[135]\, 
        \data_selected[148]\, N_672, \data_temp[103]_net_1\, 
        N_685, \data_temp[116]_net_1\, N_704, N_717, 
        \data_temp_5[71]\, \data_temp_5[84]\, \data_temp_5[103]\, 
        \data_temp_5[116]\, \data_selected[102]\, 
        \data_selected[117]\, \data_selected[134]\, 
        \data_selected[149]\, N_671, \data_temp[102]_net_1\, 
        N_686, \data_temp[117]_net_1\, N_703, N_718, 
        \data_temp_5[70]\, \data_temp_5[85]\, \data_temp_5[102]\, 
        \data_temp_5[117]\, \data_selected[101]\, 
        \data_selected[118]\, \data_selected[133]\, 
        \data_selected[150]\, N_670, \data_temp[101]_net_1\, 
        N_687, \data_temp[118]_net_1\, N_702, N_719, 
        \data_temp_5[69]\, \data_temp_5[86]\, \data_temp_5[101]\, 
        \data_temp_5[118]\, \data_selected[100]\, 
        \data_selected[119]\, \data_selected[132]\, 
        \data_selected[151]\, N_669, \data_temp[100]_net_1\, 
        N_688, \data_temp[119]_net_1\, N_701, N_720, 
        \data_temp_5[68]\, \data_temp_5[87]\, \data_temp_5[100]\, 
        \data_temp_5[119]\, \data_selected[99]\, 
        \data_selected[120]\, \data_selected[131]\, 
        \data_selected[152]\, N_668, \data_temp[99]_net_1\, N_689, 
        \data_temp[120]_net_1\, N_700, N_721, \data_temp_5[67]\, 
        \data_temp_5[88]\, \data_temp_5[99]\, \data_temp_5[120]\, 
        \data_selected[98]\, \data_selected[121]\, 
        \data_selected[130]\, \data_selected[153]\, N_667, 
        \data_temp[98]_net_1\, N_690, \data_temp[121]_net_1\, 
        N_699, N_722, \data_temp_5[66]\, \data_temp_5[89]\, 
        \data_temp_5[98]\, \data_temp_5[121]\, 
        \data_selected[97]\, \data_selected[122]\, 
        \data_selected[129]\, \data_selected[154]\, N_666, 
        \data_temp[97]_net_1\, N_691, \data_temp[122]_net_1\, 
        N_698, N_723, \data_temp_5[65]\, \data_temp_5[90]\, 
        \data_temp_5[97]\, \data_temp_5[122]\, 
        \data_selected[96]\, \data_selected[109]\, 
        \data_selected[128]\, \data_selected[141]\, N_665, 
        \data_temp[96]_net_1\, N_678, \data_temp[109]_net_1\, 
        N_697, N_710, \data_temp_5[64]\, \data_temp_5[77]\, 
        \data_temp_5[96]\, \data_temp_5[109]\, \data_wen_3[1]\, 
        \time_en_temp[1]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \data_temp_RNO_2[65]\ : MX2C
      port map(A => data_f2_out(97), B => data_f3_out(97), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_734);
    
    \data_temp[124]\ : DFN1C0
      port map(D => N_245, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[124]_net_1\);
    
    \data_temp_RNO_4[42]\ : MX2
      port map(A => data_f2_out(74), B => data_f3_out(74), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_767);
    
    \data_temp[99]\ : DFN1C0
      port map(D => \data_temp_5[99]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[99]_net_1\);
    
    \data_temp_RNO_1[76]\ : MX2C
      port map(A => N_731, B => N_806, S => N_1580_2, Y => 
        \data_selected[108]\);
    
    \data_temp_RNO_0[42]\ : AO1D
      port map(A => N_912_i, B => N_842, C => N_1668, Y => 
        \data_temp_5_i_0[42]\);
    
    \data[3]\ : DFN1C0
      port map(D => \data_5[3]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(3));
    
    \data_temp_RNO_2[32]\ : MX2
      port map(A => data_f0_out(64), B => data_f1_out(64), S => 
        \data_valid_and_ready_0[0]_net_1\, Y => N_769);
    
    \data_temp_RNO_2[64]\ : MX2C
      port map(A => data_f2_out(96), B => data_f3_out(96), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_747);
    
    \time_en_temp[1]\ : DFN1E0C0
      port map(D => N_917, CLK => HCLK_c, CLR => HRESETn_c, E => 
        state_0_sqmuxa_i, Q => \time_en_temp[1]_net_1\);
    
    \data_temp[127]\ : DFN1C0
      port map(D => \data_temp_5[127]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[127]_net_1\);
    
    \time_wen_RNO[1]\ : INV
      port map(A => N_857, Y => N_857_i);
    
    \data_RNO[13]\ : NOR2A
      port map(A => \data_temp[13]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[13]\);
    
    \state_RNIQTIC[2]\ : NOR2
      port map(A => \state[4]_net_1\, B => \state[2]_net_1\, Y
         => N_928);
    
    \data_temp_RNO_1[86]\ : MX2C
      port map(A => N_1725, B => N_802, S => N_1580_3, Y => 
        \data_selected[118]\);
    
    \data_temp_RNO_1[73]\ : MX2C
      port map(A => N_1740, B => N_817, S => N_1580_2, Y => 
        \data_selected[105]\);
    
    \data_temp_RNO_0[103]\ : MX2C
      port map(A => \data_temp[103]_net_1\, B => 
        \data_selected[135]\, S => \state[4]_net_1\, Y => N_704);
    
    \data_temp_RNO_1[101]\ : MX2C
      port map(A => N_1712, B => N_789, S => N_1580_3, Y => 
        \data_selected[133]\);
    
    \data_temp_RNO_2[124]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1693, 
        Y => N_904);
    
    \data_temp_RNO_1[96]\ : MX2C
      port map(A => N_1721, B => N_798, S => N_1580, Y => 
        \data_selected[128]\);
    
    \data_temp_RNO_1[83]\ : MX2C
      port map(A => N_1736, B => N_799, S => N_1580_3, Y => 
        \data_selected[115]\);
    
    \data_temp[26]\ : DFN1C0
      port map(D => \data_temp_5[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[26]_net_1\);
    
    \data_RNO[17]\ : NOR2A
      port map(A => \data_temp[17]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[17]\);
    
    \data_valid_ack[3]\ : DFN1E0C0
      port map(D => N_860_i, CLK => HCLK_c, CLR => HRESETn_c, E
         => N_929, Q => valid_ack(3));
    
    \data_temp_RNO_1[39]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_764, 
        Y => N_1660);
    
    \data_temp_RNO_1[93]\ : MX2
      port map(A => data_f0_out(125), B => data_f1_out(125), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_795);
    
    \data_temp[13]\ : DFN1C0
      port map(D => \data_temp_5[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[13]_net_1\);
    
    \data_temp[56]\ : DFN1C0
      port map(D => \data_temp_5[56]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[56]_net_1\);
    
    \data_temp_RNO_2[127]\ : MX2C
      port map(A => data_f2_out(159), B => data_f3_out(159), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1696);
    
    \data_temp[125]\ : DFN1C0
      port map(D => N_247, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[125]_net_1\);
    
    \data_temp_RNO[65]\ : NOR2A
      port map(A => N_863, B => N_666, Y => \data_temp_5[65]\);
    
    \data_temp_RNO[98]\ : NOR2A
      port map(A => N_863, B => N_699, Y => \data_temp_5[98]\);
    
    \data_RNO[5]\ : NOR2A
      port map(A => \data_temp[5]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[5]\);
    
    \data_temp_RNO_2[119]\ : MX2C
      port map(A => data_f2_out(151), B => data_f3_out(151), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1702);
    
    \data_wen[3]\ : DFN1E0P0
      port map(D => \data_wen_3[3]\, CLK => HCLK_c, PRE => 
        HRESETn_c, E => N_928, Q => data_wen(3));
    
    \data_temp[70]\ : DFN1C0
      port map(D => \data_temp_5[70]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[70]_net_1\);
    
    \data_temp_RNO[39]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[39]\, C => 
        N_1660, Y => N_231);
    
    \data_temp_RNO[77]\ : NOR2A
      port map(A => N_863, B => N_678, Y => \data_temp_5[77]\);
    
    \data[13]\ : DFN1C0
      port map(D => \data_5[13]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(13));
    
    \data_temp_RNO_2[57]\ : MX2C
      port map(A => data_f2_out(89), B => data_f3_out(89), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_754);
    
    \data_temp[64]\ : DFN1C0
      port map(D => \data_temp_5[64]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[64]_net_1\);
    
    \data_temp_RNO[93]\ : NOR3B
      port map(A => N_863_0, B => N_914, C => 
        \data_temp_5_i_0[93]\, Y => N_243);
    
    \state_RNO_0[4]\ : OR3
      port map(A => \state[2]_net_1\, B => \state[1]_net_1\, C
         => \state[3]_net_1\, Y => \state_ns_i_i_a2_1[0]\);
    
    \data_temp_RNO_1[50]\ : MX2C
      port map(A => N_761, B => N_836, S => N_1580_1, Y => 
        \data_selected[82]\);
    
    \data_temp[6]\ : DFN1C0
      port map(D => \data_temp_5[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[6]_net_1\);
    
    \data[31]\ : DFN1C0
      port map(D => \data_5[31]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(31));
    
    \data_temp[112]\ : DFN1C0
      port map(D => \data_temp_5[112]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[112]_net_1\);
    
    \data_temp_RNO[112]\ : NOR2A
      port map(A => N_863_1, B => N_713, Y => \data_temp_5[112]\);
    
    \data_temp[100]\ : DFN1C0
      port map(D => \data_temp_5[100]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[100]_net_1\);
    
    \data_temp_RNO_2[70]\ : MX2C
      port map(A => data_f2_out(102), B => data_f3_out(102), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_739);
    
    \data_temp_RNO_3[56]\ : MX2C
      port map(A => data_f0_out(88), B => data_f1_out(88), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_828);
    
    \data_temp_RNO_0[37]\ : AO1D
      port map(A => N_912_i, B => N_851, C => N_1653, Y => 
        \data_temp_5_i_0[37]\);
    
    \data_temp_RNO[36]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[36]\, C => 
        N_1651, Y => N_225);
    
    \data_temp_RNO_0[59]\ : MX2C
      port map(A => \data_temp[91]_net_1\, B => 
        \data_selected[91]\, S => \state[4]_net_1\, Y => N_660);
    
    \data_temp_RNO_0[51]\ : MX2C
      port map(A => \data_temp[83]_net_1\, B => 
        \data_selected[83]\, S => \state[4]_net_1\, Y => N_652);
    
    \data_temp_RNO_3[66]\ : MX2C
      port map(A => data_f0_out(98), B => data_f1_out(98), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_824);
    
    \data_temp_RNO_3[86]\ : MX2C
      port map(A => data_f0_out(118), B => data_f1_out(118), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_802);
    
    \data_temp_RNO_3[49]\ : MX2C
      port map(A => data_f0_out(81), B => data_f1_out(81), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_835);
    
    \data_temp_RNO_3[41]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[73]_net_1\, 
        Y => N_1665);
    
    \data_temp_RNO_2[40]\ : MX2
      port map(A => data_f0_out(72), B => data_f1_out(72), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_854);
    
    \data_temp_RNO_0[116]\ : MX2C
      port map(A => \data_temp[116]_net_1\, B => 
        \data_selected[148]\, S => \state[4]_net_1\, Y => N_717);
    
    \data_temp_RNO_1[35]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1688, 
        Y => N_874);
    
    \data_temp_RNO_3[53]\ : MX2C
      port map(A => data_f0_out(85), B => data_f1_out(85), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_839);
    
    \data_temp_RNO[49]\ : NOR2A
      port map(A => N_863_1, B => N_650, Y => \data_temp_5[49]\);
    
    \data_temp_RNO_3[63]\ : MX2C
      port map(A => data_f0_out(95), B => data_f1_out(95), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_821);
    
    \data_temp_RNO_3[83]\ : MX2C
      port map(A => data_f0_out(115), B => data_f1_out(115), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_799);
    
    \data_temp_RNO_2[120]\ : MX2C
      port map(A => data_f2_out(152), B => data_f3_out(152), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1703);
    
    \data_temp_RNO_1[52]\ : MX2C
      port map(A => N_749, B => N_838, S => N_1580_1, Y => 
        \data_selected[84]\);
    
    \data_temp_RNO_1[34]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1687, 
        Y => N_871);
    
    \state[2]\ : DFN1C0
      port map(D => \state[3]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[2]_net_1\);
    
    \data_temp[36]\ : DFN1C0
      port map(D => N_225, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[36]_net_1\);
    
    un5_data_selected_i_i_a2 : OR2B
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_917);
    
    \data_wen_RNO[0]\ : OR2
      port map(A => \time_en_temp[0]_net_1\, B => 
        \state[4]_net_1\, Y => \data_wen_3[0]\);
    
    \data_temp_RNO_2[72]\ : MX2C
      port map(A => data_f2_out(104), B => data_f3_out(104), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1739);
    
    \data_temp_RNO_1[110]\ : MX2C
      port map(A => N_1707, B => N_784, S => N_1580_2, Y => 
        \data_selected[142]\);
    
    \data_temp[82]\ : DFN1C0
      port map(D => \data_temp_5[82]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[82]_net_1\);
    
    \data_temp_RNO[46]\ : NOR2A
      port map(A => N_863_0, B => N_647, Y => \data_temp_5[46]\);
    
    \data_temp[0]\ : DFN1C0
      port map(D => \data_temp_5[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[0]_net_1\);
    
    data_selected_sn_m2_0_o2_2 : OR2A
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_1580_2);
    
    \data_temp_RNO_2[42]\ : MX2
      port map(A => data_f0_out(74), B => data_f1_out(74), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_842);
    
    \data_temp_RNO_1[49]\ : MX2C
      port map(A => N_760, B => N_835, S => N_1580_1, Y => 
        \data_selected[81]\);
    
    \data_temp_RNO_1[41]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_766, 
        Y => N_1666);
    
    \data_RNO[2]\ : NOR2A
      port map(A => \data_temp[2]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[2]\);
    
    \data_temp_RNO_2[86]\ : MX2C
      port map(A => data_f2_out(118), B => data_f3_out(118), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1725);
    
    \data_temp[10]\ : DFN1C0
      port map(D => \data_temp_5[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[10]_net_1\);
    
    \data_temp[111]\ : DFN1C0
      port map(D => \data_temp_5[111]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[111]_net_1\);
    
    \data_temp_RNO_3[36]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[68]_net_1\, 
        Y => N_1650);
    
    \data_temp_RNO_0[55]\ : MX2C
      port map(A => \data_temp[87]_net_1\, B => 
        \data_selected[87]\, S => \state[4]_net_1\, Y => N_656);
    
    \time_wen[1]\ : DFN1E0P0
      port map(D => N_857_i, CLK => HCLK_c, PRE => HRESETn_c, E
         => N_928, Q => time_wen(1));
    
    \data_temp_RNO_1[127]\ : MX2C
      port map(A => N_1696, B => N_1684, S => N_1580_1, Y => 
        \data_selected[159]\);
    
    \data_temp_RNO[10]\ : NOR2A
      port map(A => \data_temp[42]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[10]\);
    
    \data_temp_RNO_3[45]\ : MX2C
      port map(A => data_f0_out(77), B => data_f1_out(77), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_845);
    
    \data_temp_RNO_3[108]\ : MX2C
      port map(A => data_f0_out(140), B => data_f1_out(140), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_782);
    
    \data_temp[24]\ : DFN1C0
      port map(D => \data_temp_5[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[24]_net_1\);
    
    \data_temp_RNO_0[115]\ : MX2C
      port map(A => \data_temp[115]_net_1\, B => 
        \data_selected[147]\, S => \state[4]_net_1\, Y => N_716);
    
    \data_temp_RNO_2[83]\ : MX2C
      port map(A => data_f2_out(115), B => data_f3_out(115), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1736);
    
    \data_temp_RNO_0[54]\ : MX2C
      port map(A => \data_temp[86]_net_1\, B => 
        \data_selected[86]\, S => \state[4]_net_1\, Y => N_655);
    
    \data_temp_RNO[4]\ : NOR2A
      port map(A => \data_temp[36]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[4]\);
    
    \data_temp[119]\ : DFN1C0
      port map(D => \data_temp_5[119]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[119]_net_1\);
    
    \data_temp_RNO_3[33]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[65]_net_1\, 
        Y => N_867);
    
    \data_temp_RNO_2[66]\ : MX2C
      port map(A => data_f2_out(98), B => data_f3_out(98), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_735);
    
    \data_temp[54]\ : DFN1C0
      port map(D => \data_temp_5[54]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[54]_net_1\);
    
    \data_temp_RNO_3[44]\ : MX2C
      port map(A => data_f0_out(76), B => data_f1_out(76), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_844);
    
    \data_temp_RNO[75]\ : NOR2A
      port map(A => N_863_2, B => N_676, Y => \data_temp_5[75]\);
    
    \data_temp[81]\ : DFN1C0
      port map(D => \data_temp_5[81]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[81]_net_1\);
    
    \data_RNO[11]\ : NOR2A
      port map(A => \data_temp[11]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[11]\);
    
    \data_temp_RNO_3[99]\ : MX2C
      port map(A => data_f0_out(131), B => data_f1_out(131), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_787);
    
    \data_temp_RNO_3[91]\ : MX2
      port map(A => data_f2_out(123), B => data_f3_out(123), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1730);
    
    \data_temp_RNO[37]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[37]\, C => 
        N_1654, Y => N_227);
    
    \data_temp_RNO_2[63]\ : MX2C
      port map(A => data_f2_out(95), B => data_f3_out(95), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_746);
    
    \data_RNO[12]\ : NOR2A
      port map(A => \data_temp[12]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[12]\);
    
    \data_valid_ack_RNO[0]\ : INV
      port map(A => \time_wen_3[0]\, Y => \time_wen_3_i[0]\);
    
    \data_temp_RNO_3[127]\ : MX2C
      port map(A => data_f0_out(159), B => data_f1_out(159), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1684);
    
    \data_temp_RNO[2]\ : NOR2A
      port map(A => \data_temp[34]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[2]\);
    
    \data_temp_RNO_1[68]\ : MX2C
      port map(A => N_737, B => N_826, S => N_1580_3, Y => 
        \data_selected[100]\);
    
    \data_temp_RNO_0[120]\ : MX2C
      port map(A => \data_temp[120]_net_1\, B => 
        \data_selected[152]\, S => \state[4]_net_1\, Y => N_721);
    
    \data_temp_RNO_1[45]\ : MX2C
      port map(A => N_756, B => N_845, S => N_1580_1, Y => 
        \data_selected[77]\);
    
    \data_temp_RNO_0[98]\ : MX2C
      port map(A => \data_temp[98]_net_1\, B => 
        \data_selected[130]\, S => \state[4]_net_1\, Y => N_699);
    
    \data_temp_RNO[91]\ : NOR3B
      port map(A => N_863_0, B => N_913, C => 
        \data_temp_5_i_0[91]\, Y => N_249);
    
    \data_temp_RNO[115]\ : NOR2A
      port map(A => N_863_2, B => N_716, Y => \data_temp_5[115]\);
    
    \data_temp[76]\ : DFN1C0
      port map(D => \data_temp_5[76]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[76]_net_1\);
    
    \data_temp_RNO_1[44]\ : MX2C
      port map(A => N_755, B => N_844, S => N_1580_1, Y => 
        \data_selected[76]\);
    
    \data_RNO[28]\ : NOR2A
      port map(A => \data_temp[28]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[28]\);
    
    \data_temp_RNO[68]\ : NOR2A
      port map(A => N_863, B => N_669, Y => \data_temp_5[68]\);
    
    \data_temp_RNO_0[117]\ : MX2C
      port map(A => \data_temp[117]_net_1\, B => 
        \data_selected[149]\, S => \state[4]_net_1\, Y => N_718);
    
    \data_temp_RNO[92]\ : NOR3B
      port map(A => N_863_0, B => N_915, C => 
        \data_temp_5_i_0[92]\, Y => N_241);
    
    \time_en_temp_RNO[2]\ : OR2
      port map(A => \data_valid_and_ready_0[2]_net_1\, B => 
        N_1580_0, Y => N_858);
    
    \data_temp_RNO_3[122]\ : MX2C
      port map(A => data_f0_out(154), B => data_f1_out(154), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1679);
    
    \data_temp_RNO_2[50]\ : MX2C
      port map(A => data_f2_out(82), B => data_f3_out(82), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_761);
    
    \data_temp[88]\ : DFN1C0
      port map(D => \data_temp_5[88]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[88]_net_1\);
    
    \data[28]\ : DFN1C0
      port map(D => \data_5[28]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(28));
    
    \data_temp_RNO[20]\ : NOR2A
      port map(A => \data_temp[52]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[20]\);
    
    \data_temp_RNO[63]\ : NOR2A
      port map(A => N_863_1, B => N_664, Y => \data_temp_5[63]\);
    
    \data_temp_RNO[47]\ : NOR2A
      port map(A => N_863_0, B => N_648, Y => \data_temp_5[47]\);
    
    \data_temp_RNO[117]\ : NOR2A
      port map(A => N_863_2, B => N_718, Y => \data_temp_5[117]\);
    
    \data_wen_RNO[1]\ : OR2
      port map(A => \time_en_temp[1]_net_1\, B => 
        \state[4]_net_1\, Y => \data_wen_3[1]\);
    
    \data_temp[93]\ : DFN1C0
      port map(D => N_243, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[93]_net_1\);
    
    \data_temp[49]\ : DFN1C0
      port map(D => \data_temp_5[49]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[49]_net_1\);
    
    \data_temp_RNO_3[95]\ : MX2C
      port map(A => data_f0_out(127), B => data_f1_out(127), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_797);
    
    \data_temp_RNO_2[109]\ : MX2C
      port map(A => data_f2_out(141), B => data_f3_out(141), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1706);
    
    \data[5]\ : DFN1C0
      port map(D => \data_5[5]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(5));
    
    \data_temp_RNO_4[41]\ : MX2
      port map(A => data_f2_out(73), B => data_f3_out(73), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_766);
    
    \data_temp[34]\ : DFN1C0
      port map(D => N_221, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[34]_net_1\);
    
    \data[16]\ : DFN1C0
      port map(D => \data_5[16]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(16));
    
    \data_temp_RNO_3[78]\ : MX2C
      port map(A => data_f0_out(110), B => data_f1_out(110), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_808);
    
    \data_temp_RNO_0[49]\ : MX2C
      port map(A => \data_temp[81]_net_1\, B => 
        \data_selected[81]\, S => \state[4]_net_1\, Y => N_650);
    
    \data_temp_RNO_0[41]\ : AO1D
      port map(A => N_912_i, B => N_841, C => N_1665, Y => 
        \data_temp_5_i_0[41]\);
    
    \data_temp[62]\ : DFN1C0
      port map(D => \data_temp_5[62]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[62]_net_1\);
    
    \data_temp_RNO[94]\ : NOR2A
      port map(A => N_863_1, B => N_695, Y => \data_temp_5[94]\);
    
    \data[7]\ : DFN1C0
      port map(D => \data_5[7]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(7));
    
    \data_temp_RNO_3[114]\ : MX2C
      port map(A => data_f0_out(146), B => data_f1_out(146), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_774);
    
    \data_temp_RNO_2[39]\ : MX2
      port map(A => data_f0_out(71), B => data_f1_out(71), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_853);
    
    \data_temp_RNO[122]\ : NOR2A
      port map(A => N_863, B => N_723, Y => \data_temp_5[122]\);
    
    \data_RNO[31]\ : NOR2A
      port map(A => \data_temp[31]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[31]\);
    
    \data_temp_RNO_3[94]\ : MX2C
      port map(A => data_f0_out(126), B => data_f1_out(126), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_796);
    
    \data_temp[87]\ : DFN1C0
      port map(D => \data_temp_5[87]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[87]_net_1\);
    
    \data_temp_RNO_3[126]\ : MX2C
      port map(A => data_f0_out(158), B => data_f1_out(158), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1683);
    
    \data_temp_RNO_0[78]\ : MX2C
      port map(A => \data_temp[110]_net_1\, B => 
        \data_selected[110]\, S => \state[4]_net_1\, Y => N_679);
    
    \data_temp_RNO_2[52]\ : MX2C
      port map(A => data_f2_out(84), B => data_f3_out(84), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_749);
    
    \data_temp[108]\ : DFN1C0
      port map(D => \data_temp_5[108]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[108]_net_1\);
    
    \data_temp_RNO_1[112]\ : MX2C
      port map(A => N_1709, B => N_772, S => N_1580_2, Y => 
        \data_selected[144]\);
    
    \data_temp_RNO_0[106]\ : MX2C
      port map(A => \data_temp[106]_net_1\, B => 
        \data_selected[138]\, S => \state[4]_net_1\, Y => N_707);
    
    \data_temp_RNO[59]\ : NOR2A
      port map(A => N_863_1, B => N_660, Y => \data_temp_5[59]\);
    
    \data_temp_RNO_0[32]\ : AO1D
      port map(A => N_912_i, B => N_769, C => N_864, Y => 
        \data_temp_5_i_0[32]\);
    
    \data_temp[61]\ : DFN1C0
      port map(D => \data_temp_5[61]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[61]_net_1\);
    
    \data_temp_RNO_4[38]\ : MX2
      port map(A => data_f2_out(70), B => data_f3_out(70), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_763);
    
    \data_temp[16]\ : DFN1C0
      port map(D => \data_temp_5[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[16]_net_1\);
    
    \data[21]\ : DFN1C0
      port map(D => \data_5[21]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(21));
    
    \data_temp_RNO_1[36]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1689, 
        Y => N_1651);
    
    \data_temp_RNO[89]\ : NOR2A
      port map(A => N_863, B => N_690, Y => \data_temp_5[89]\);
    
    \data_temp_RNO[35]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[35]\, C => 
        N_874, Y => N_223);
    
    \data_temp_RNO[102]\ : NOR2A
      port map(A => N_863_2, B => N_703, Y => \data_temp_5[102]\);
    
    \data_temp_RNO_1[123]\ : MX2
      port map(A => data_f0_out(155), B => data_f1_out(155), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1680);
    
    \data_temp_RNO_3[110]\ : MX2C
      port map(A => data_f0_out(142), B => data_f1_out(142), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_784);
    
    \data_temp_RNO_2[122]\ : MX2C
      port map(A => data_f2_out(154), B => data_f3_out(154), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1691);
    
    \data_temp_RNO_0[45]\ : MX2C
      port map(A => \data_temp[77]_net_1\, B => 
        \data_selected[77]\, S => \state[4]_net_1\, Y => N_646);
    
    \data_temp_RNO_2[125]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1694, 
        Y => N_906);
    
    \data[0]\ : DFN1C0
      port map(D => \data_5[0]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(0));
    
    \data_temp_RNO[56]\ : NOR2A
      port map(A => N_863_1, B => N_657, Y => \data_temp_5[56]\);
    
    \data_temp_RNO_2[35]\ : MX2
      port map(A => data_f0_out(67), B => data_f1_out(67), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_849);
    
    \data_valid_ack[0]\ : DFN1E0C0
      port map(D => \time_wen_3_i[0]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_929, Q => valid_ack(0));
    
    \data_temp_RNO_1[33]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1686, 
        Y => N_868);
    
    \data_temp_RNO[86]\ : NOR2A
      port map(A => N_863, B => N_687, Y => \data_temp_5[86]\);
    
    \data_temp_RNO_1[119]\ : MX2C
      port map(A => N_1702, B => N_1676, S => N_1580, Y => 
        \data_selected[151]\);
    
    \data_temp_RNO_1[100]\ : MX2C
      port map(A => N_1711, B => N_788, S => N_1580, Y => 
        \data_selected[132]\);
    
    \data_temp_RNO_1[118]\ : MX2C
      port map(A => N_1701, B => N_1675, S => N_1580_3, Y => 
        \data_selected[150]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \data_temp_RNO_0[44]\ : MX2C
      port map(A => \data_temp[76]_net_1\, B => 
        \data_selected[76]\, S => \state[4]_net_1\, Y => N_645);
    
    \data_temp_RNO_2[34]\ : MX2
      port map(A => data_f0_out(66), B => data_f1_out(66), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_848);
    
    \data_RNO[16]\ : NOR2A
      port map(A => \data_temp[16]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[16]\);
    
    \data_temp[74]\ : DFN1C0
      port map(D => \data_temp_5[74]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[74]_net_1\);
    
    \data_temp[90]\ : DFN1C0
      port map(D => \data_temp_5[90]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[90]_net_1\);
    
    \data_temp[22]\ : DFN1C0
      port map(D => \data_temp_5[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[22]_net_1\);
    
    \time_wen_3_i_a2_0[3]\ : NOR2B
      port map(A => \data_valid_and_ready[3]_net_1\, B => 
        \data_valid_and_ready_0[2]_net_1\, Y => 
        \time_wen_3_i_a2_0[3]_net_1\);
    
    \state_RNIUI96[4]\ : CLKINT
      port map(A => \state_0[4]\, Y => \state[4]_net_1\);
    
    \data_temp_RNO_0[56]\ : MX2C
      port map(A => \data_temp[88]_net_1\, B => 
        \data_selected[88]\, S => \state[4]_net_1\, Y => N_657);
    
    \data_temp_RNO_0[88]\ : MX2C
      port map(A => \data_temp[120]_net_1\, B => 
        \data_selected[120]\, S => \state[4]_net_1\, Y => N_689);
    
    \data_temp_RNO[78]\ : NOR2A
      port map(A => N_863_1, B => N_679, Y => \data_temp_5[78]\);
    
    \data_temp_RNO_1[67]\ : MX2C
      port map(A => N_736, B => N_825, S => N_1580, Y => 
        \data_selected[99]\);
    
    \data_temp_RNO[45]\ : NOR2A
      port map(A => N_863_0, B => N_646, Y => \data_temp_5[45]\);
    
    \data_temp_RNO_3[46]\ : MX2C
      port map(A => data_f0_out(78), B => data_f1_out(78), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_846);
    
    \data_temp_RNO_0[112]\ : MX2C
      port map(A => \data_temp[112]_net_1\, B => 
        \data_selected[144]\, S => \state[4]_net_1\, Y => N_713);
    
    \data_temp[68]\ : DFN1C0
      port map(D => \data_temp_5[68]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[68]_net_1\);
    
    \time_en_temp[2]\ : DFN1E0C0
      port map(D => N_858, CLK => HCLK_c, CLR => HRESETn_c, E => 
        state_0_sqmuxa_i, Q => \time_en_temp[2]_net_1\);
    
    \data_temp_RNO_2[98]\ : MX2C
      port map(A => data_f2_out(130), B => data_f3_out(130), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1723);
    
    \data_temp_RNO_0[105]\ : MX2C
      port map(A => \data_temp[105]_net_1\, B => 
        \data_selected[137]\, S => \state[4]_net_1\, Y => N_706);
    
    \data_temp_RNIDNBC[124]\ : OR2
      port map(A => \state[4]_net_1\, B => \data_temp[124]_net_1\, 
        Y => N_915);
    
    \data_temp[52]\ : DFN1C0
      port map(D => \data_temp_5[52]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[52]_net_1\);
    
    \data_temp_RNO_0[97]\ : MX2C
      port map(A => \data_temp[97]_net_1\, B => 
        \data_selected[129]\, S => \state[4]_net_1\, Y => N_698);
    
    \data_temp_RNO_0[119]\ : MX2C
      port map(A => \data_temp[119]_net_1\, B => 
        \data_selected[151]\, S => \state[4]_net_1\, Y => N_720);
    
    \data[2]\ : DFN1C0
      port map(D => \data_5[2]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(2));
    
    \data_temp_RNO[73]\ : NOR2A
      port map(A => N_863_2, B => N_674, Y => \data_temp_5[73]\);
    
    \data_temp[85]\ : DFN1C0
      port map(D => \data_temp_5[85]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[85]_net_1\);
    
    \data_temp_5_i_a2_0_0[32]\ : NOR2A
      port map(A => \data_valid_and_ready_0[2]_net_1\, B => 
        \data_valid_and_ready[3]_net_1\, Y => 
        \data_temp_5_i_a2_0_0[32]_net_1\);
    
    \data_valid_and_ready_1[2]\ : OR2A
      port map(A => valid_out_2, B => ready_i_0(2), Y => 
        \data_valid_and_ready_1[2]_net_1\);
    
    \data_temp_RNO_0[53]\ : MX2C
      port map(A => \data_temp[85]_net_1\, B => 
        \data_selected[85]\, S => \state[4]_net_1\, Y => N_654);
    
    \data_temp_RNO_3[43]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[75]_net_1\, 
        Y => N_897);
    
    \data[22]\ : DFN1C0
      port map(D => \data_5[22]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(22));
    
    \data_temp_RNO_2[126]\ : MX2C
      port map(A => data_f2_out(158), B => data_f3_out(158), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1695);
    
    \data_temp_RNO[61]\ : NOR2A
      port map(A => N_863_1, B => N_662, Y => \data_temp_5[61]\);
    
    \data_temp_RNO_0[68]\ : MX2C
      port map(A => \data_temp[100]_net_1\, B => 
        \data_selected[100]\, S => \state[4]_net_1\, Y => N_669);
    
    \data_temp[67]\ : DFN1C0
      port map(D => \data_temp_5[67]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[67]_net_1\);
    
    \data_temp[21]\ : DFN1C0
      port map(D => \data_temp_5[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[21]_net_1\);
    
    \data_wen[2]\ : DFN1E0P0
      port map(D => \data_wen_3[2]\, CLK => HCLK_c, PRE => 
        HRESETn_c, E => N_928, Q => data_wen(2));
    
    \data_temp[9]\ : DFN1C0
      port map(D => \data_temp_5[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[9]_net_1\);
    
    \data_temp_RNO[62]\ : NOR2A
      port map(A => N_863_1, B => N_663, Y => \data_temp_5[62]\);
    
    \data_temp_RNO[125]\ : NOR3B
      port map(A => N_863_0, B => N_914, C => 
        \data_temp_5_i_0[125]\, Y => N_247);
    
    \data_temp_RNO_1[59]\ : MX2C
      port map(A => N_742, B => N_831, S => N_1580_2, Y => 
        \data_selected[91]\);
    
    \data_temp_RNO_1[51]\ : MX2C
      port map(A => N_748, B => N_837, S => N_1580_1, Y => 
        \data_selected[83]\);
    
    \data_temp_RNO_1[46]\ : MX2C
      port map(A => N_757, B => N_846, S => N_1580_1, Y => 
        \data_selected[78]\);
    
    \data_temp[51]\ : DFN1C0
      port map(D => \data_temp_5[51]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[51]_net_1\);
    
    data_selected_sn_m2_0_o2_3 : OR2A
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_1580_3);
    
    \data_temp_RNO_2[79]\ : MX2C
      port map(A => data_f2_out(111), B => data_f3_out(111), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1732);
    
    \data_temp_RNO_2[71]\ : MX2C
      port map(A => data_f2_out(103), B => data_f3_out(103), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_740);
    
    \data_temp_RNO_3[77]\ : MX2C
      port map(A => data_f0_out(109), B => data_f1_out(109), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_807);
    
    \data_temp[120]\ : DFN1C0
      port map(D => \data_temp_5[120]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[120]_net_1\);
    
    \state_RNIKK3V21_3[4]\ : OR3B
      port map(A => \state[4]_net_1\, B => 
        \time_wen_3_i_a2_0[3]_net_1\, C => N_1580_0, Y => N_860);
    
    \data_temp[106]\ : DFN1C0
      port map(D => \data_temp_5[106]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[106]_net_1\);
    
    \time_wen[3]\ : DFN1E0P0
      port map(D => N_860, CLK => HCLK_c, PRE => HRESETn_c, E => 
        N_928, Q => time_wen(3));
    
    \data_temp_RNO_2[49]\ : MX2C
      port map(A => data_f2_out(81), B => data_f3_out(81), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_760);
    
    \data_temp_RNO_2[41]\ : MX2
      port map(A => data_f0_out(73), B => data_f1_out(73), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_841);
    
    \data_temp_RNO[127]\ : NOR2A
      port map(A => N_863_0, B => N_728, Y => \data_temp_5[127]\);
    
    \data_temp_RNO_0[107]\ : MX2C
      port map(A => \data_temp[107]_net_1\, B => 
        \data_selected[139]\, S => \state[4]_net_1\, Y => N_708);
    
    \data_temp_RNO_0[77]\ : MX2C
      port map(A => \data_temp[109]_net_1\, B => 
        \data_selected[109]\, S => \state[4]_net_1\, Y => N_678);
    
    \data_temp_RNO_1[43]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_768, 
        Y => N_898);
    
    \data_temp_RNO[57]\ : NOR2A
      port map(A => N_863_1, B => N_658, Y => \data_temp_5[57]\);
    
    \data_temp_RNO[64]\ : NOR2A
      port map(A => N_863, B => N_665, Y => \data_temp_5[64]\);
    
    \data_temp[14]\ : DFN1C0
      port map(D => \data_temp_5[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[14]_net_1\);
    
    \data_temp_RNO[87]\ : NOR2A
      port map(A => N_863, B => N_688, Y => \data_temp_5[87]\);
    
    \data_temp[114]\ : DFN1C0
      port map(D => \data_temp_5[114]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[114]_net_1\);
    
    \data_temp_RNO_0[124]\ : AO1D
      port map(A => N_1681, B => N_912_i, C => N_904, Y => 
        \data_temp_5_i_0[124]\);
    
    \data_temp_RNO[110]\ : NOR2A
      port map(A => N_863_1, B => N_711, Y => \data_temp_5[110]\);
    
    \data_temp_RNO_3[111]\ : MX2C
      port map(A => data_f0_out(143), B => data_f1_out(143), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_771);
    
    \data_temp_RNO_0[121]\ : MX2C
      port map(A => \data_temp[121]_net_1\, B => 
        \data_selected[153]\, S => \state[4]_net_1\, Y => N_722);
    
    \data_temp_RNO[105]\ : NOR2A
      port map(A => N_863_2, B => N_706, Y => \data_temp_5[105]\);
    
    \data[29]\ : DFN1C0
      port map(D => \data_5[29]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(29));
    
    \data_temp_RNO_1[78]\ : MX2C
      port map(A => N_733, B => N_808, S => N_1580_2, Y => 
        \data_selected[110]\);
    
    \data_temp[32]\ : DFN1C0
      port map(D => N_215, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[32]_net_1\);
    
    \data_temp_RNO_0[118]\ : MX2C
      port map(A => \data_temp[118]_net_1\, B => 
        \data_selected[150]\, S => \state[4]_net_1\, Y => N_719);
    
    \data_temp[28]\ : DFN1C0
      port map(D => \data_temp_5[28]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[28]_net_1\);
    
    \data_temp_RNO_3[96]\ : MX2C
      port map(A => data_f0_out(128), B => data_f1_out(128), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_798);
    
    \data_temp[117]\ : DFN1C0
      port map(D => \data_temp_5[117]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[117]_net_1\);
    
    \data_RNO[19]\ : NOR2A
      port map(A => \data_temp[19]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[19]\);
    
    \data_temp_RNO_4[37]\ : MX2
      port map(A => data_f2_out(69), B => data_f3_out(69), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_762);
    
    data_selected_sn_m2_0_o2 : OR2A
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_1580);
    
    \data_temp[58]\ : DFN1C0
      port map(D => \data_temp_5[58]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[58]_net_1\);
    
    \data_temp_RNO_1[55]\ : MX2C
      port map(A => N_752, B => N_827, S => N_1580_1, Y => 
        \data_selected[87]\);
    
    \data_temp_RNO_3[104]\ : MX2C
      port map(A => data_f0_out(136), B => data_f1_out(136), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_778);
    
    \data_temp_RNO_1[88]\ : MX2C
      port map(A => N_1727, B => N_804, S => N_1580, Y => 
        \data_selected[120]\);
    
    \data_temp_RNO[107]\ : NOR2A
      port map(A => N_863_2, B => N_708, Y => \data_temp_5[107]\);
    
    \state_RNIKK3V21_1[4]\ : OR3B
      port map(A => \state[4]_net_1\, B => 
        \data_temp_5_i_a2_0_0[32]_net_1\, C => N_1580_0, Y => 
        N_863_2);
    
    \data[25]\ : DFN1C0
      port map(D => \data_5[25]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(25));
    
    \data_temp_RNO_3[93]\ : MX2
      port map(A => data_f2_out(125), B => data_f3_out(125), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1718);
    
    \data_temp_RNO_2[75]\ : MX2C
      port map(A => data_f2_out(107), B => data_f3_out(107), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_730);
    
    \data_valid_and_ready_0[2]\ : OR2A
      port map(A => valid_out_2, B => ready_i_0(2), Y => 
        \data_valid_and_ready_0[2]_net_1\);
    
    \data_temp_RNO_1[115]\ : MX2C
      port map(A => N_1698, B => N_775, S => N_1580_3, Y => 
        \data_selected[147]\);
    
    \data_temp[27]\ : DFN1C0
      port map(D => \data_temp_5[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[27]_net_1\);
    
    \data_temp_RNO_1[54]\ : MX2C
      port map(A => N_751, B => N_840, S => N_1580_1, Y => 
        \data_selected[86]\);
    
    \data_temp_RNO[38]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[38]\, C => 
        N_1657, Y => N_229);
    
    \data_temp_RNO_2[45]\ : MX2C
      port map(A => data_f2_out(77), B => data_f3_out(77), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_756);
    
    \data_temp_RNO_1[98]\ : MX2C
      port map(A => N_1723, B => N_786, S => N_1580, Y => 
        \data_selected[130]\);
    
    \data_temp[31]\ : DFN1C0
      port map(D => \data_temp_5[31]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[31]_net_1\);
    
    \data_temp_RNO_1[102]\ : MX2C
      port map(A => N_1713, B => N_790, S => N_1580_3, Y => 
        \data_selected[134]\);
    
    \data_temp[3]\ : DFN1C0
      port map(D => \data_temp_5[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[3]_net_1\);
    
    \data_temp_RNO_2[74]\ : MX2C
      port map(A => data_f2_out(106), B => data_f3_out(106), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_729);
    
    \data_temp[65]\ : DFN1C0
      port map(D => \data_temp_5[65]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[65]_net_1\);
    
    \data_temp[57]\ : DFN1C0
      port map(D => \data_temp_5[57]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[57]_net_1\);
    
    \state_RNIHQ76Q[4]\ : OR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_859);
    
    \data_temp_RNO_3[115]\ : MX2C
      port map(A => data_f0_out(147), B => data_f1_out(147), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_775);
    
    \state_RNO[3]\ : INV
      port map(A => state_0_sqmuxa_i, Y => state_0_sqmuxa_i_i);
    
    \data_temp[7]\ : DFN1C0
      port map(D => \data_temp_5[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[7]_net_1\);
    
    \data_temp_RNO[33]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[33]\, C => 
        N_868, Y => N_219);
    
    \data_temp_RNO_2[44]\ : MX2C
      port map(A => data_f2_out(76), B => data_f3_out(76), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_755);
    
    \data_temp_RNO_2[118]\ : MX2C
      port map(A => data_f2_out(150), B => data_f3_out(150), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1701);
    
    \data_temp_RNO_1[116]\ : MX2C
      port map(A => N_1699, B => N_776, S => N_1580_3, Y => 
        \data_selected[148]\);
    
    \data_temp[96]\ : DFN1C0
      port map(D => \data_temp_5[96]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[96]_net_1\);
    
    \data_temp_RNO_0[87]\ : MX2C
      port map(A => \data_temp[119]_net_1\, B => 
        \data_selected[119]\, S => \state[4]_net_1\, Y => N_688);
    
    \data_temp[115]\ : DFN1C0
      port map(D => \data_temp_5[115]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[115]_net_1\);
    
    \data_temp_RNO_3[100]\ : MX2C
      port map(A => data_f0_out(132), B => data_f1_out(132), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_788);
    
    \data[14]\ : DFN1C0
      port map(D => \data_5[14]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(14));
    
    \data_temp_RNO_2[97]\ : MX2C
      port map(A => data_f2_out(129), B => data_f3_out(129), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1722);
    
    \data_temp_RNO_0[123]\ : AO1D
      port map(A => N_1680, B => N_912_i, C => N_910, Y => 
        \data_temp_5_i_0[123]\);
    
    \data_temp_RNO[71]\ : NOR2A
      port map(A => N_863_2, B => N_672, Y => \data_temp_5[71]\);
    
    \data_temp[43]\ : DFN1C0
      port map(D => N_239, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[43]_net_1\);
    
    \data_temp_RNO_0[46]\ : MX2C
      port map(A => \data_temp[78]_net_1\, B => 
        \data_selected[78]\, S => \state[4]_net_1\, Y => N_647);
    
    \data_temp_RNO_1[60]\ : MX2C
      port map(A => N_743, B => N_832, S => N_1580_2, Y => 
        \data_selected[92]\);
    
    \data_temp_RNO_1[121]\ : MX2C
      port map(A => N_1690, B => N_1678, S => N_1580, Y => 
        \data_selected[153]\);
    
    \data_temp_RNO_2[36]\ : MX2
      port map(A => data_f0_out(68), B => data_f1_out(68), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_850);
    
    \data_temp_RNO[72]\ : NOR2A
      port map(A => N_863_2, B => N_673, Y => \data_temp_5[72]\);
    
    \data_temp_RNO[116]\ : NOR2A
      port map(A => N_863_2, B => N_717, Y => \data_temp_5[116]\);
    
    \data_temp_RNO_0[90]\ : MX2C
      port map(A => \data_temp[122]_net_1\, B => 
        \data_selected[122]\, S => \state[4]_net_1\, Y => N_691);
    
    \data_RNO[24]\ : NOR2A
      port map(A => \data_temp[24]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[24]\);
    
    \data_temp_RNO_1[109]\ : MX2C
      port map(A => N_1706, B => N_783, S => N_1580, Y => 
        \data_selected[141]\);
    
    \data_temp_RNO[90]\ : NOR2A
      port map(A => N_863, B => N_691, Y => \data_temp_5[90]\);
    
    \data_temp_RNO[48]\ : NOR2A
      port map(A => N_863_1, B => N_649, Y => \data_temp_5[48]\);
    
    \data_temp_RNO_1[108]\ : MX2C
      port map(A => N_1705, B => N_782, S => N_1580_2, Y => 
        \data_selected[140]\);
    
    \data_temp[72]\ : DFN1C0
      port map(D => \data_temp_5[72]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[72]_net_1\);
    
    \data_temp_RNO_2[111]\ : MX2C
      port map(A => data_f2_out(143), B => data_f3_out(143), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1708);
    
    \data_temp_RNO[5]\ : NOR2A
      port map(A => \data_temp[37]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[5]\);
    
    \data_temp_RNO_4[43]\ : MX2
      port map(A => data_f2_out(75), B => data_f3_out(75), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_768);
    
    \data_temp_RNO[55]\ : NOR2A
      port map(A => N_863_1, B => N_656, Y => \data_temp_5[55]\);
    
    \data_temp_RNO_0[67]\ : MX2C
      port map(A => \data_temp[99]_net_1\, B => 
        \data_selected[99]\, S => \state[4]_net_1\, Y => N_668);
    
    \data_temp_RNO_0[43]\ : AO1D
      port map(A => N_912_i, B => N_843, C => N_897, Y => 
        \data_temp_5_i_0[43]\);
    
    \data_temp[38]\ : DFN1C0
      port map(D => N_229, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[38]_net_1\);
    
    \data_RNO[20]\ : NOR2A
      port map(A => \data_temp[20]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[20]\);
    
    \data_temp_RNO[85]\ : NOR2A
      port map(A => N_863_2, B => N_686, Y => \data_temp_5[85]\);
    
    \data_temp_RNO[7]\ : NOR2A
      port map(A => \data_temp[39]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[7]\);
    
    \data_temp_RNO[43]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[43]\, C => 
        N_898, Y => N_239);
    
    \data_temp[103]\ : DFN1C0
      port map(D => \data_temp_5[103]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[103]_net_1\);
    
    \data[10]\ : DFN1C0
      port map(D => \data_5[10]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(10));
    
    \data_temp_RNO_2[33]\ : MX2
      port map(A => data_f0_out(65), B => data_f1_out(65), S => 
        \data_valid_and_ready_0[0]_net_1\, Y => N_770);
    
    \data_temp_RNO_3[58]\ : MX2C
      port map(A => data_f0_out(90), B => data_f1_out(90), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_830);
    
    \data_temp_RNO_3[68]\ : MX2C
      port map(A => data_f0_out(100), B => data_f1_out(100), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_826);
    
    \data_temp_RNO_0[102]\ : MX2C
      port map(A => \data_temp[102]_net_1\, B => 
        \data_selected[134]\, S => \state[4]_net_1\, Y => N_703);
    
    \state[4]\ : DFN1P0
      port map(D => N_861, CLK => HCLK_c, PRE => HRESETn_c, Q => 
        \state_0[4]\);
    
    \data_temp_RNO_3[88]\ : MX2C
      port map(A => data_f0_out(120), B => data_f1_out(120), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_804);
    
    \data_temp_RNO[74]\ : NOR2A
      port map(A => N_863_2, B => N_675, Y => \data_temp_5[74]\);
    
    \data_temp_RNO_2[59]\ : MX2C
      port map(A => data_f2_out(91), B => data_f3_out(91), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_742);
    
    \data_temp_RNO_2[51]\ : MX2C
      port map(A => data_f2_out(83), B => data_f3_out(83), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_748);
    
    \data_temp_RNO_0[109]\ : MX2C
      port map(A => \data_temp[109]_net_1\, B => 
        \data_selected[141]\, S => \state[4]_net_1\, Y => N_710);
    
    \data_temp_RNO_3[113]\ : MX2C
      port map(A => data_f0_out(145), B => data_f1_out(145), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_773);
    
    \data_temp_RNO_1[62]\ : MX2C
      port map(A => N_745, B => N_820, S => N_1580_2, Y => 
        \data_selected[94]\);
    
    \data_temp_RNO_1[114]\ : MX2C
      port map(A => N_1697, B => N_774, S => N_1580_3, Y => 
        \data_selected[146]\);
    
    \data_temp_RNO_0[92]\ : AO1D
      port map(A => N_912_i, B => N_794, C => N_900, Y => 
        \data_temp_5_i_0[92]\);
    
    \data_valid_and_ready[3]\ : NOR2B
      port map(A => valid_out_3, B => ready_i_0(3), Y => 
        \data_valid_and_ready[3]_net_1\);
    
    \data_temp[37]\ : DFN1C0
      port map(D => N_227, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[37]_net_1\);
    
    \data_temp[71]\ : DFN1C0
      port map(D => \data_temp_5[71]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[71]_net_1\);
    
    \data_temp_RNO_3[70]\ : MX2C
      port map(A => data_f0_out(102), B => data_f1_out(102), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_814);
    
    \data_temp_RNO_0[39]\ : AO1D
      port map(A => N_912_i, B => N_853, C => N_1659, Y => 
        \data_temp_5_i_0[39]\);
    
    \state_RNIR1JC[3]\ : NOR2
      port map(A => \state[4]_net_1\, B => \state[3]_net_1\, Y
         => N_929);
    
    \data_temp[25]\ : DFN1C0
      port map(D => \data_temp_5[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[25]_net_1\);
    
    \data_temp_RNO[9]\ : NOR2A
      port map(A => \data_temp[41]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[9]\);
    
    \data_RNO[25]\ : NOR2A
      port map(A => \data_temp[25]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[25]\);
    
    \data_temp_RNO_0[70]\ : MX2C
      port map(A => \data_temp[102]_net_1\, B => 
        \data_selected[102]\, S => \state[4]_net_1\, Y => N_671);
    
    \data_temp[55]\ : DFN1C0
      port map(D => \data_temp_5[55]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[55]_net_1\);
    
    \data_temp_RNO_1[77]\ : MX2C
      port map(A => N_732, B => N_807, S => N_1580, Y => 
        \data_selected[109]\);
    
    \data_temp_RNO_2[88]\ : MX2C
      port map(A => data_f2_out(120), B => data_f3_out(120), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1727);
    
    \data_temp_RNO_2[113]\ : MX2C
      port map(A => data_f2_out(145), B => data_f3_out(145), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1710);
    
    \data_temp_RNO_3[38]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[70]_net_1\, 
        Y => N_1656);
    
    \data_temp[40]\ : DFN1C0
      port map(D => N_233, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[40]_net_1\);
    
    \data_temp_RNO[120]\ : NOR2A
      port map(A => N_863, B => N_721, Y => \data_temp_5[120]\);
    
    \data_temp_RNO_1[87]\ : MX2C
      port map(A => N_1726, B => N_803, S => N_1580_3, Y => 
        \data_selected[119]\);
    
    \data_temp[12]\ : DFN1C0
      port map(D => \data_temp_5[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[12]_net_1\);
    
    \data_temp_RNO_2[55]\ : MX2C
      port map(A => data_f2_out(87), B => data_f3_out(87), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_752);
    
    \data_temp_RNO_3[72]\ : MX2C
      port map(A => data_f0_out(104), B => data_f1_out(104), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_816);
    
    \data_wen[1]\ : DFN1E0P0
      port map(D => \data_wen_3[1]\, CLK => HCLK_c, PRE => 
        HRESETn_c, E => N_928, Q => data_wen(1));
    
    \data_temp_RNO[19]\ : NOR2A
      port map(A => \data_temp[51]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[19]\);
    
    \data_temp[94]\ : DFN1C0
      port map(D => \data_temp_5[94]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[94]_net_1\);
    
    \data_temp[78]\ : DFN1C0
      port map(D => \data_temp_5[78]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[78]_net_1\);
    
    \data_temp_RNO_2[68]\ : MX2C
      port map(A => data_f2_out(100), B => data_f3_out(100), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_737);
    
    \data_temp_RNO_3[101]\ : MX2C
      port map(A => data_f0_out(133), B => data_f1_out(133), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_789);
    
    \data_temp_RNO_2[54]\ : MX2C
      port map(A => data_f2_out(86), B => data_f3_out(86), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_751);
    
    \data_temp_RNO_1[97]\ : MX2C
      port map(A => N_1722, B => N_785, S => N_1580, Y => 
        \data_selected[129]\);
    
    \data_temp_RNO_0[72]\ : MX2C
      port map(A => \data_temp[104]_net_1\, B => 
        \data_selected[104]\, S => \state[4]_net_1\, Y => N_673);
    
    \data_temp_RNO_0[35]\ : AO1D
      port map(A => N_912_i, B => N_849, C => N_873, Y => 
        \data_temp_5_i_0[35]\);
    
    \data_RNO[7]\ : NOR2A
      port map(A => \data_temp[7]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[7]\);
    
    \data_temp_RNO[31]\ : NOR2A
      port map(A => \data_temp[63]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[31]\);
    
    \data_temp_RNO_0[108]\ : MX2C
      port map(A => \data_temp[108]_net_1\, B => 
        \data_selected[140]\, S => \state[4]_net_1\, Y => N_709);
    
    \data[27]\ : DFN1C0
      port map(D => \data_5[27]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(27));
    
    \data_temp_RNICJBC[123]\ : OR2
      port map(A => \state[4]_net_1\, B => \data_temp[123]_net_1\, 
        Y => N_913);
    
    \data_temp[5]\ : DFN1C0
      port map(D => \data_temp_5[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[5]_net_1\);
    
    \data_temp_RNO[32]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[32]\, C => 
        N_865, Y => N_215);
    
    \data_temp_RNO[16]\ : NOR2A
      port map(A => \data_temp[48]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[16]\);
    
    \data_temp_RNO_0[34]\ : AO1D
      port map(A => N_912_i, B => N_848, C => N_870, Y => 
        \data_temp_5_i_0[34]\);
    
    \data_temp_RNO[100]\ : NOR2A
      port map(A => N_863, B => N_701, Y => \data_temp_5[100]\);
    
    \state[1]\ : DFN1C0
      port map(D => \state[2]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[1]_net_1\);
    
    \data_temp[102]\ : DFN1C0
      port map(D => \data_temp_5[102]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[102]_net_1\);
    
    \data_temp_RNO_1[56]\ : MX2C
      port map(A => N_753, B => N_828, S => N_1580_1, Y => 
        \data_selected[88]\);
    
    \data_temp[77]\ : DFN1C0
      port map(D => \data_temp_5[77]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[77]_net_1\);
    
    \data_temp[11]\ : DFN1C0
      port map(D => \data_temp_5[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[11]_net_1\);
    
    \data_temp[89]\ : DFN1C0
      port map(D => \data_temp_5[89]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[89]_net_1\);
    
    \data_RNO[0]\ : NOR2A
      port map(A => \data_temp[0]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[0]\);
    
    \data_temp_RNO_4[32]\ : MX2
      port map(A => data_f2_out(64), B => data_f3_out(64), S => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_1685);
    
    \data_temp_RNO[118]\ : NOR2A
      port map(A => N_863, B => N_719, Y => \data_temp_5[118]\);
    
    \data_temp_RNO_2[76]\ : MX2C
      port map(A => data_f2_out(108), B => data_f3_out(108), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_731);
    
    \data_temp_RNO_0[80]\ : MX2C
      port map(A => \data_temp[112]_net_1\, B => 
        \data_selected[112]\, S => \state[4]_net_1\, Y => N_681);
    
    \data_temp_RNO_1[105]\ : MX2C
      port map(A => N_1716, B => N_779, S => N_1580_3, Y => 
        \data_selected[137]\);
    
    \data_temp[35]\ : DFN1C0
      port map(D => N_223, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[35]_net_1\);
    
    \data_temp_RNO_2[90]\ : MX2C
      port map(A => data_f2_out(122), B => data_f3_out(122), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1729);
    
    \data_temp_RNO_2[114]\ : MX2C
      port map(A => data_f2_out(146), B => data_f3_out(146), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1697);
    
    data_selected_sn_m2_0_o2_1 : OR2A
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_1580_1);
    
    \data_temp_RNO_2[46]\ : MX2C
      port map(A => data_f2_out(78), B => data_f3_out(78), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_757);
    
    \data_valid_and_ready_2[0]\ : OR2A
      port map(A => valid_out_0, B => ready_i_0(0), Y => 
        \data_valid_and_ready_2[0]_net_1\);
    
    \data_temp_RNO_1[53]\ : MX2C
      port map(A => N_750, B => N_839, S => N_1580_1, Y => 
        \data_selected[85]\);
    
    \data_temp_RNO[34]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[34]\, C => 
        N_871, Y => N_221);
    
    \data_temp_RNO[0]\ : NOR2A
      port map(A => \data_temp[32]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[0]\);
    
    \data_temp_RNO[41]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[41]\, C => 
        N_1666, Y => N_235);
    
    \data_temp_RNO_3[105]\ : MX2C
      port map(A => data_f0_out(137), B => data_f1_out(137), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_779);
    
    \data[8]\ : DFN1C0
      port map(D => \data_5[8]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(8));
    
    \data_temp_RNO_2[73]\ : MX2C
      port map(A => data_f2_out(105), B => data_f3_out(105), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1740);
    
    state_0_sqmuxa_i_0_o2_0_a2 : NOR2
      port map(A => \data_valid_and_ready[3]_net_1\, B => N_916, 
        Y => N_1306);
    
    \data_temp_RNO_2[108]\ : MX2C
      port map(A => data_f2_out(140), B => data_f3_out(140), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1705);
    
    \data_temp_RNO[60]\ : NOR2A
      port map(A => N_863_1, B => N_661, Y => \data_temp_5[60]\);
    
    \data_temp_RNO_1[106]\ : MX2C
      port map(A => N_1717, B => N_780, S => N_1580_2, Y => 
        \data_selected[138]\);
    
    \data_temp_RNO[42]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[42]\, C => 
        N_1669, Y => N_237);
    
    \data_temp_RNO_2[43]\ : MX2
      port map(A => data_f0_out(75), B => data_f1_out(75), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_843);
    
    \data_RNO[4]\ : NOR2A
      port map(A => \data_temp[4]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[4]\);
    
    \data_temp_RNO_3[57]\ : MX2C
      port map(A => data_f0_out(89), B => data_f1_out(89), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_829);
    
    \data_temp_RNO[126]\ : NOR2A
      port map(A => N_863_1, B => N_727, Y => \data_temp_5[126]\);
    
    \data_temp_RNO_0[60]\ : MX2C
      port map(A => \data_temp[92]_net_1\, B => 
        \data_selected[92]\, S => \state[4]_net_1\, Y => N_661);
    
    \data_temp_RNO_3[67]\ : MX2C
      port map(A => data_f0_out(99), B => data_f1_out(99), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_825);
    
    \data_temp_RNO_2[117]\ : MX2C
      port map(A => data_f2_out(149), B => data_f3_out(149), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1700);
    
    \data_temp_RNO_3[87]\ : MX2C
      port map(A => data_f0_out(119), B => data_f1_out(119), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_803);
    
    \data_temp_RNO[58]\ : NOR2A
      port map(A => N_863_1, B => N_659, Y => \data_temp_5[58]\);
    
    \data_temp[2]\ : DFN1C0
      port map(D => \data_temp_5[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[2]_net_1\);
    
    \data_temp_RNO[29]\ : NOR2A
      port map(A => \data_temp[61]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[29]\);
    
    \data_temp[18]\ : DFN1C0
      port map(D => \data_temp_5[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[18]_net_1\);
    
    \data_temp_RNO_0[82]\ : MX2C
      port map(A => \data_temp[114]_net_1\, B => 
        \data_selected[114]\, S => \state[4]_net_1\, Y => N_683);
    
    \data_temp_RNO[88]\ : NOR2A
      port map(A => N_863, B => N_689, Y => \data_temp_5[88]\);
    
    \data_temp_RNO_2[92]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1731, 
        Y => N_900);
    
    \data_temp_RNO[8]\ : NOR2A
      port map(A => \data_temp[40]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[8]\);
    
    \data_temp[101]\ : DFN1C0
      port map(D => \data_temp_5[101]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[101]_net_1\);
    
    \data_temp_RNO_2[101]\ : MX2C
      port map(A => data_f2_out(133), B => data_f3_out(133), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1712);
    
    \data_temp_RNO[53]\ : NOR2A
      port map(A => N_863_1, B => N_654, Y => \data_temp_5[53]\);
    
    \data_temp_RNO[44]\ : NOR2A
      port map(A => N_863_0, B => N_645, Y => \data_temp_5[44]\);
    
    \data_temp_RNO[83]\ : NOR2A
      port map(A => N_863_2, B => N_684, Y => \data_temp_5[83]\);
    
    \time_en_temp[0]\ : DFN1E0C0
      port map(D => \data_valid_and_ready[0]_net_1\, CLK => 
        HCLK_c, CLR => HRESETn_c, E => state_0_sqmuxa_i, Q => 
        \time_en_temp[0]_net_1\);
    
    \data_temp_RNO[26]\ : NOR2A
      port map(A => \data_temp[58]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[26]\);
    
    \data_temp[126]\ : DFN1C0
      port map(D => \data_temp_5[126]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[126]_net_1\);
    
    \data_temp_RNO[106]\ : NOR2A
      port map(A => N_863_2, B => N_707, Y => \data_temp_5[106]\);
    
    \data_temp[17]\ : DFN1C0
      port map(D => \data_temp_5[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[17]_net_1\);
    
    \data_temp[109]\ : DFN1C0
      port map(D => \data_temp_5[109]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[109]_net_1\);
    
    \data_temp_RNO_0[62]\ : MX2C
      port map(A => \data_temp[94]_net_1\, B => 
        \data_selected[94]\, S => \state[4]_net_1\, Y => N_663);
    
    \data_RNO[23]\ : NOR2A
      port map(A => \data_temp[23]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[23]\);
    
    \data[6]\ : DFN1C0
      port map(D => \data_5[6]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(6));
    
    \data_temp_RNO[17]\ : NOR2A
      port map(A => \data_temp[49]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[17]\);
    
    un23_data_selected_i_a2 : OR2A
      port map(A => \data_valid_and_ready_0[2]_net_1\, B => 
        N_1580_1, Y => N_916);
    
    \data_temp_RNO_2[87]\ : MX2C
      port map(A => data_f2_out(119), B => data_f3_out(119), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1726);
    
    \data_temp_RNO[114]\ : NOR2A
      port map(A => N_863_2, B => N_715, Y => \data_temp_5[114]\);
    
    \data_temp_RNO_3[103]\ : MX2C
      port map(A => data_f0_out(135), B => data_f1_out(135), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_791);
    
    \data_temp_RNO_1[70]\ : MX2C
      port map(A => N_739, B => N_814, S => N_1580_3, Y => 
        \data_selected[102]\);
    
    \data_temp[75]\ : DFN1C0
      port map(D => \data_temp_5[75]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[75]_net_1\);
    
    \data_temp_RNO_3[37]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[69]_net_1\, 
        Y => N_1653);
    
    \data_temp_RNO_1[38]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_763, 
        Y => N_1657);
    
    \data_temp_RNO_1[104]\ : MX2C
      port map(A => N_1715, B => N_778, S => N_1580_3, Y => 
        \data_selected[136]\);
    
    \state_RNIKK3V21_0[4]\ : OR3B
      port map(A => \state[4]_net_1\, B => 
        \data_temp_5_i_a2_0_0[32]_net_1\, C => N_1580_0, Y => 
        N_863_1);
    
    \data_temp[46]\ : DFN1C0
      port map(D => \data_temp_5[46]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[46]_net_1\);
    
    \data_temp_RNO[111]\ : NOR2A
      port map(A => N_863_2, B => N_712, Y => \data_temp_5[111]\);
    
    \data_temp_RNO_2[110]\ : MX2C
      port map(A => data_f2_out(142), B => data_f3_out(142), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1707);
    
    \data_temp[69]\ : DFN1C0
      port map(D => \data_temp_5[69]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[69]_net_1\);
    
    \data_temp_RNO_1[80]\ : MX2C
      port map(A => N_1733, B => N_810, S => N_1580_2, Y => 
        \data_selected[112]\);
    
    \data_temp_RNO_2[67]\ : MX2C
      port map(A => data_f2_out(99), B => data_f3_out(99), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_736);
    
    \data_RNO[27]\ : NOR2A
      port map(A => \data_temp[27]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[27]\);
    
    \data_temp_RNO[6]\ : NOR2A
      port map(A => \data_temp[38]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[6]\);
    
    \data_temp_RNO_0[126]\ : MX2C
      port map(A => \data_temp[126]_net_1\, B => 
        \data_selected[158]\, S => \state[4]_net_1\, Y => N_727);
    
    \data_temp_RNO_1[90]\ : MX2C
      port map(A => N_1729, B => N_792, S => N_1580, Y => 
        \data_selected[122]\);
    
    \data[23]\ : DFN1C0
      port map(D => \data_5[23]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(23));
    
    \data_temp_RNO_2[103]\ : MX2C
      port map(A => data_f2_out(135), B => data_f3_out(135), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1714);
    
    \state_RNIKK3V21[4]\ : OR3B
      port map(A => \state[4]_net_1\, B => 
        \data_temp_5_i_a2_0_0[32]_net_1\, C => N_1580_0, Y => 
        N_863_0);
    
    \data_temp_RNO_1[72]\ : MX2C
      port map(A => N_1739, B => N_816, S => N_1580_3, Y => 
        \data_selected[104]\);
    
    \data_temp_RNO_0[58]\ : MX2C
      port map(A => \data_temp[90]_net_1\, B => 
        \data_selected[90]\, S => \state[4]_net_1\, Y => N_659);
    
    \data_temp_RNO_1[117]\ : MX2C
      port map(A => N_1700, B => N_777, S => N_1580_3, Y => 
        \data_selected[149]\);
    
    \data_temp[4]\ : DFN1C0
      port map(D => \data_temp_5[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[4]_net_1\);
    
    \data_wen_RNO[2]\ : OR2
      port map(A => \time_en_temp[2]_net_1\, B => 
        \state[4]_net_1\, Y => \data_wen_3[2]\);
    
    \data_temp_RNO_3[48]\ : MX2C
      port map(A => data_f0_out(80), B => data_f1_out(80), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_834);
    
    \data_temp[92]\ : DFN1C0
      port map(D => N_241, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[92]_net_1\);
    
    \data_temp_RNO_2[56]\ : MX2C
      port map(A => data_f2_out(88), B => data_f3_out(88), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_753);
    
    \state_RNIKK3V21_2[4]\ : OR3B
      port map(A => \state[4]_net_1\, B => 
        \data_temp_5_i_a2_0_0[32]_net_1\, C => N_1580_0, Y => 
        N_863);
    
    \data_temp_RNO[70]\ : NOR2A
      port map(A => N_863_2, B => N_671, Y => \data_temp_5[70]\);
    
    \data_temp_RNO_1[82]\ : MX2C
      port map(A => N_1735, B => N_812, S => N_1580_3, Y => 
        \data_selected[114]\);
    
    \data_RNO[18]\ : NOR2A
      port map(A => \data_temp[18]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[18]\);
    
    \time_wen[0]\ : DFN1E0P0
      port map(D => \time_wen_3[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, E => N_928, Q => time_wen(0));
    
    \data_temp_RNO_1[120]\ : MX2C
      port map(A => N_1703, B => N_1677, S => N_1580, Y => 
        \data_selected[152]\);
    
    \data_temp_RNO_0[36]\ : AO1D
      port map(A => N_912_i, B => N_850, C => N_1650, Y => 
        \data_temp_5_i_0[36]\);
    
    \data_temp_RNO_2[53]\ : MX2C
      port map(A => data_f2_out(85), B => data_f3_out(85), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_750);
    
    \data_temp_RNO_1[69]\ : MX2C
      port map(A => N_738, B => N_813, S => N_1580_3, Y => 
        \data_selected[101]\);
    
    \data_temp_RNO_1[61]\ : MX2C
      port map(A => N_744, B => N_833, S => N_1580_2, Y => 
        \data_selected[93]\);
    
    \state[0]\ : DFN1C0
      port map(D => \state[1]_net_1\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[0]_net_1\);
    
    \data_temp_RNO[27]\ : NOR2A
      port map(A => \data_temp[59]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[27]\);
    
    \data_temp_RNO_1[92]\ : MX2
      port map(A => data_f0_out(124), B => data_f1_out(124), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_794);
    
    \data_temp_RNO_0[99]\ : MX2C
      port map(A => \data_temp[99]_net_1\, B => 
        \data_selected[131]\, S => \state[4]_net_1\, Y => N_700);
    
    \data_temp_RNO_0[91]\ : AO1D
      port map(A => N_912_i, B => N_793, C => N_908, Y => 
        \data_temp_5_i_0[91]\);
    
    \data_temp[15]\ : DFN1C0
      port map(D => \data_temp_5[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[15]_net_1\);
    
    \data_temp_RNO[119]\ : NOR2A
      port map(A => N_863, B => N_720, Y => \data_temp_5[119]\);
    
    \data_RNO[1]\ : NOR2A
      port map(A => \data_temp[1]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[1]\);
    
    \data_temp_RNO_3[117]\ : MX2C
      port map(A => data_f0_out(149), B => data_f1_out(149), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_777);
    
    \data_temp_RNO_0[33]\ : AO1D
      port map(A => N_912_i, B => N_770, C => N_867, Y => 
        \data_temp_5_i_0[33]\);
    
    \data_temp[91]\ : DFN1C0
      port map(D => N_249, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[91]_net_1\);
    
    \data_temp_RNO_0[125]\ : AO1D
      port map(A => N_1682, B => N_912_i, C => N_906, Y => 
        \data_temp_5_i_0[125]\);
    
    \data_temp_RNO_0[110]\ : MX2C
      port map(A => \data_temp[110]_net_1\, B => 
        \data_selected[142]\, S => \state[4]_net_1\, Y => N_711);
    
    \data_temp_RNO_1[48]\ : MX2C
      port map(A => N_759, B => N_834, S => N_1580_1, Y => 
        \data_selected[80]\);
    
    \data_temp_RNO[15]\ : NOR2A
      port map(A => \data_temp[47]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[15]\);
    
    \data[18]\ : DFN1C0
      port map(D => \data_5[18]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(18));
    
    \data_temp[29]\ : DFN1C0
      port map(D => \data_temp_5[29]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[29]_net_1\);
    
    \data_temp_RNO_3[50]\ : MX2C
      port map(A => data_f0_out(82), B => data_f1_out(82), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_836);
    
    \data_temp[110]\ : DFN1C0
      port map(D => \data_temp_5[110]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[110]_net_1\);
    
    data_selected_sn_m2_0_o2_0 : OR2A
      port map(A => \data_valid_and_ready_0[0]_net_1\, B => 
        \data_valid_and_ready[1]_net_1\, Y => N_1580_0);
    
    \data_temp_RNO[51]\ : NOR2A
      port map(A => N_863_1, B => N_652, Y => \data_temp_5[51]\);
    
    \data_temp_RNO[113]\ : NOR2A
      port map(A => N_863_2, B => N_714, Y => \data_temp_5[113]\);
    
    \data_temp_RNO_3[60]\ : MX2C
      port map(A => data_f0_out(92), B => data_f1_out(92), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_832);
    
    \data_temp[123]\ : DFN1C0
      port map(D => N_251, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[123]_net_1\);
    
    \data_temp_RNO_3[80]\ : MX2C
      port map(A => data_f0_out(112), B => data_f1_out(112), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_810);
    
    \data_temp_RNO_2[104]\ : MX2C
      port map(A => data_f2_out(136), B => data_f3_out(136), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1715);
    
    \data_temp_RNO[81]\ : NOR2A
      port map(A => N_863_2, B => N_682, Y => \data_temp_5[81]\);
    
    \data_temp_RNO[1]\ : NOR2A
      port map(A => \data_temp[33]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[1]\);
    
    \data_temp[59]\ : DFN1C0
      port map(D => \data_temp_5[59]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[59]_net_1\);
    
    \data_temp_RNO[52]\ : NOR2A
      port map(A => N_863_1, B => N_653, Y => \data_temp_5[52]\);
    
    \data_temp_RNO[82]\ : NOR2A
      port map(A => N_863_2, B => N_683, Y => \data_temp_5[82]\);
    
    \data_temp_RNO[108]\ : NOR2A
      port map(A => N_863_1, B => N_709, Y => \data_temp_5[108]\);
    
    \data_temp_RNO_3[112]\ : MX2C
      port map(A => data_f0_out(144), B => data_f1_out(144), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_772);
    
    \data_temp_RNO_3[79]\ : MX2C
      port map(A => data_f0_out(111), B => data_f1_out(111), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_809);
    
    \data_temp_RNO_3[71]\ : MX2C
      port map(A => data_f0_out(103), B => data_f1_out(103), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_815);
    
    \data_temp[44]\ : DFN1C0
      port map(D => \data_temp_5[44]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[44]_net_1\);
    
    \data_temp_RNO_1[65]\ : MX2C
      port map(A => N_734, B => N_823, S => N_1580, Y => 
        \data_selected[97]\);
    
    \data_temp_RNO_2[107]\ : MX2C
      port map(A => data_f2_out(139), B => data_f3_out(139), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1704);
    
    \data_temp_RNO_3[98]\ : MX2C
      port map(A => data_f0_out(130), B => data_f1_out(130), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_786);
    
    \data_temp_RNO_0[95]\ : MX2C
      port map(A => \data_temp[127]_net_1\, B => 
        \data_selected[127]\, S => \state[4]_net_1\, Y => N_696);
    
    \data_temp_RNO_0[79]\ : MX2C
      port map(A => \data_temp[111]_net_1\, B => 
        \data_selected[111]\, S => \state[4]_net_1\, Y => N_680);
    
    \data_temp_RNO_0[71]\ : MX2C
      port map(A => \data_temp[103]_net_1\, B => 
        \data_selected[103]\, S => \state[4]_net_1\, Y => N_672);
    
    \data_valid_ack_RNO[3]\ : INV
      port map(A => N_860, Y => N_860_i);
    
    \data_temp_RNO_3[52]\ : MX2C
      port map(A => data_f0_out(84), B => data_f1_out(84), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_838);
    
    \data_temp[98]\ : DFN1C0
      port map(D => \data_temp_5[98]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[98]_net_1\);
    
    \data_temp_RNO[54]\ : NOR2A
      port map(A => N_863_1, B => N_655, Y => \data_temp_5[54]\);
    
    \data_valid_and_ready_1[0]\ : OR2A
      port map(A => valid_out_0, B => ready_i_0(0), Y => 
        \data_valid_and_ready_1[0]_net_1\);
    
    \data_temp_RNO_3[62]\ : MX2C
      port map(A => data_f0_out(94), B => data_f1_out(94), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_820);
    
    \data_temp_RNO_1[37]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_762, 
        Y => N_1654);
    
    \data_temp_RNO_3[82]\ : MX2C
      port map(A => data_f0_out(114), B => data_f1_out(114), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_812);
    
    \data_temp_RNO_1[64]\ : MX2C
      port map(A => N_747, B => N_822, S => N_1580, Y => 
        \data_selected[96]\);
    
    \data_temp_RNO[84]\ : NOR2A
      port map(A => N_863_2, B => N_685, Y => \data_temp_5[84]\);
    
    \data_temp_RNO_2[80]\ : MX2C
      port map(A => data_f2_out(112), B => data_f3_out(112), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1733);
    
    \data_temp_RNO_0[94]\ : MX2C
      port map(A => \data_temp[126]_net_1\, B => 
        \data_selected[126]\, S => \state[4]_net_1\, Y => N_695);
    
    \data_temp_RNO_0[127]\ : MX2C
      port map(A => \data_temp[127]_net_1\, B => 
        \data_selected[159]\, S => \state[4]_net_1\, Y => N_728);
    
    \data_temp[83]\ : DFN1C0
      port map(D => \data_temp_5[83]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[83]_net_1\);
    
    \data_temp_RNO_3[116]\ : MX2C
      port map(A => data_f0_out(148), B => data_f1_out(148), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_776);
    
    \data[4]\ : DFN1C0
      port map(D => \data_5[4]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(4));
    
    \data[11]\ : DFN1C0
      port map(D => \data_5[11]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(11));
    
    \data_temp_RNO[124]\ : NOR3B
      port map(A => N_863_0, B => N_915, C => 
        \data_temp_5_i_0[124]\, Y => N_245);
    
    \data_valid_and_ready_3[0]\ : OR2A
      port map(A => valid_out_0, B => ready_i_0(0), Y => 
        \data_valid_and_ready_3[0]_net_1\);
    
    \data_RNO[21]\ : NOR2A
      port map(A => \data_temp[21]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[21]\);
    
    \data_temp_RNO_4[39]\ : MX2
      port map(A => data_f2_out(71), B => data_f3_out(71), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_764);
    
    \data_temp[97]\ : DFN1C0
      port map(D => \data_temp_5[97]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[97]_net_1\);
    
    \state_RNIKK3V21_4[4]\ : OR2A
      port map(A => \state[4]_net_1\, B => N_1306, Y => 
        state_0_sqmuxa_i);
    
    \data_RNO[22]\ : NOR2A
      port map(A => \data_temp[22]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[22]\);
    
    \data_temp_RNO_2[60]\ : MX2C
      port map(A => data_f2_out(92), B => data_f3_out(92), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_743);
    
    \data_temp_RNO[30]\ : NOR2A
      port map(A => \data_temp[62]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[30]\);
    
    \data_temp_RNO[25]\ : NOR2A
      port map(A => \data_temp[57]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[25]\);
    
    \data_temp_RNO[121]\ : NOR2A
      port map(A => N_863, B => N_722, Y => \data_temp_5[121]\);
    
    \time_en_temp[3]\ : DFN1E0C0
      port map(D => N_916, CLK => HCLK_c, CLR => HRESETn_c, E => 
        state_0_sqmuxa_i, Q => \time_en_temp[3]_net_1\);
    
    \data_temp_RNO_3[75]\ : MX2C
      port map(A => data_f0_out(107), B => data_f1_out(107), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_819);
    
    \data_temp_RNO_3[124]\ : MX2
      port map(A => data_f2_out(156), B => data_f3_out(156), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1693);
    
    \data_temp_RNO_0[57]\ : MX2C
      port map(A => \data_temp[89]_net_1\, B => 
        \data_selected[89]\, S => \state[4]_net_1\, Y => N_658);
    
    \data_temp[39]\ : DFN1C0
      port map(D => N_231, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[39]_net_1\);
    
    \data_temp_RNO_3[47]\ : MX2C
      port map(A => data_f0_out(79), B => data_f1_out(79), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_847);
    
    \data_temp_RNO_1[113]\ : MX2C
      port map(A => N_1710, B => N_773, S => N_1580_2, Y => 
        \data_selected[145]\);
    
    \data_temp_RNO_2[82]\ : MX2C
      port map(A => data_f2_out(114), B => data_f3_out(114), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1735);
    
    \data_temp_RNO_0[75]\ : MX2C
      port map(A => \data_temp[107]_net_1\, B => 
        \data_selected[107]\, S => \state[4]_net_1\, Y => N_676);
    
    \data_temp_RNO_3[32]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[64]_net_1\, 
        Y => N_864);
    
    \data_temp_RNO_3[74]\ : MX2C
      port map(A => data_f0_out(106), B => data_f1_out(106), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_818);
    
    \data_temp_RNO_2[100]\ : MX2C
      port map(A => data_f2_out(132), B => data_f3_out(132), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1711);
    
    \data_temp_RNO_2[112]\ : MX2C
      port map(A => data_f2_out(144), B => data_f3_out(144), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1709);
    
    \data_temp_RNO_0[48]\ : MX2C
      port map(A => \data_temp[80]_net_1\, B => 
        \data_selected[80]\, S => \state[4]_net_1\, Y => N_649);
    
    \data_temp_RNO_2[115]\ : MX2C
      port map(A => data_f2_out(147), B => data_f3_out(147), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1698);
    
    \data_temp_RNO[104]\ : NOR2A
      port map(A => N_863_2, B => N_705, Y => \data_temp_5[104]\);
    
    \data_temp_RNO_2[38]\ : MX2
      port map(A => data_f0_out(70), B => data_f1_out(70), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_852);
    
    \data_temp[122]\ : DFN1C0
      port map(D => \data_temp_5[122]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[122]_net_1\);
    
    \data_temp[8]\ : DFN1C0
      port map(D => \data_temp_5[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[8]_net_1\);
    
    \data[26]\ : DFN1C0
      port map(D => \data_5[26]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(26));
    
    \data_temp_RNO_0[74]\ : MX2C
      port map(A => \data_temp[106]_net_1\, B => 
        \data_selected[106]\, S => \state[4]_net_1\, Y => N_675);
    
    \data_temp_RNO_1[122]\ : MX2C
      port map(A => N_1691, B => N_1679, S => N_1580, Y => 
        \data_selected[154]\);
    
    \data_temp_RNO_0[89]\ : MX2C
      port map(A => \data_temp[121]_net_1\, B => 
        \data_selected[121]\, S => \state[4]_net_1\, Y => N_690);
    
    \data_temp_RNO_0[81]\ : MX2C
      port map(A => \data_temp[113]_net_1\, B => 
        \data_selected[113]\, S => \state[4]_net_1\, Y => N_682);
    
    \data_temp_RNO[101]\ : NOR2A
      port map(A => N_863, B => N_702, Y => \data_temp_5[101]\);
    
    \data_temp_RNO_2[99]\ : MX2C
      port map(A => data_f2_out(131), B => data_f3_out(131), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1724);
    
    \data_temp_RNO_2[91]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1730, 
        Y => N_908);
    
    \data_temp_RNO_2[62]\ : MX2C
      port map(A => data_f2_out(94), B => data_f3_out(94), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_745);
    
    \data_temp_RNO_3[119]\ : MX2C
      port map(A => data_f0_out(151), B => data_f1_out(151), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1676);
    
    \data_temp_RNO[40]\ : NOR3A
      port map(A => N_863_0, B => \data_temp_5_i_0[40]\, C => 
        N_1663, Y => N_233);
    
    \data_temp_RNO[99]\ : NOR2A
      port map(A => N_863, B => N_700, Y => \data_temp_5[99]\);
    
    \data_temp_RNO_4[35]\ : MX2
      port map(A => data_f2_out(67), B => data_f3_out(67), S => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_1688);
    
    \data[12]\ : DFN1C0
      port map(D => \data_5[12]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(12));
    
    \data_temp_RNO_1[107]\ : MX2C
      port map(A => N_1704, B => N_781, S => N_1580_2, Y => 
        \data_selected[139]\);
    
    \data_temp[104]\ : DFN1C0
      port map(D => \data_temp_5[104]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[104]_net_1\);
    
    \data_temp_RNO_3[120]\ : MX2C
      port map(A => data_f0_out(152), B => data_f1_out(152), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1677);
    
    \data_temp_RNO_1[47]\ : MX2C
      port map(A => N_758, B => N_847, S => N_1580_1, Y => 
        \data_selected[79]\);
    
    \data_temp_RNO_4[34]\ : MX2
      port map(A => data_f2_out(66), B => data_f3_out(66), S => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_1687);
    
    \data_temp_RNO_0[69]\ : MX2C
      port map(A => \data_temp[101]_net_1\, B => 
        \data_selected[101]\, S => \state[4]_net_1\, Y => N_670);
    
    \data_temp_RNO_0[61]\ : MX2C
      port map(A => \data_temp[93]_net_1\, B => 
        \data_selected[93]\, S => \state[4]_net_1\, Y => N_662);
    
    \data_temp_RNO[96]\ : NOR2A
      port map(A => N_863, B => N_697, Y => \data_temp_5[96]\);
    
    \data_temp[107]\ : DFN1C0
      port map(D => \data_temp_5[107]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[107]_net_1\);
    
    \data_temp[80]\ : DFN1C0
      port map(D => \data_temp_5[80]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[80]_net_1\);
    
    \data_temp_RNO_2[116]\ : MX2C
      port map(A => data_f2_out(148), B => data_f3_out(148), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1699);
    
    \data_temp_RNO[18]\ : NOR2A
      port map(A => \data_temp[50]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[18]\);
    
    \data_temp[95]\ : DFN1C0
      port map(D => \data_temp_5[95]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[95]_net_1\);
    
    \data_temp[63]\ : DFN1C0
      port map(D => \data_temp_5[63]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[63]_net_1\);
    
    \state_RNI8220I[4]\ : OR2B
      port map(A => \state[4]_net_1\, B => N_1580_1, Y => N_912_i);
    
    \data_temp_RNO[123]\ : NOR3B
      port map(A => N_863_0, B => N_913, C => 
        \data_temp_5_i_0[123]\, Y => N_251);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \data_temp_RNO_0[85]\ : MX2C
      port map(A => \data_temp[117]_net_1\, B => 
        \data_selected[117]\, S => \state[4]_net_1\, Y => N_686);
    
    \data_temp[121]\ : DFN1C0
      port map(D => \data_temp_5[121]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[121]_net_1\);
    
    \data_temp[79]\ : DFN1C0
      port map(D => \data_temp_5[79]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[79]_net_1\);
    
    \data_temp_RNO_3[107]\ : MX2C
      port map(A => data_f0_out(139), B => data_f1_out(139), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_781);
    
    \data[30]\ : DFN1C0
      port map(D => \data_5[30]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(30));
    
    \data_temp_RNO_0[122]\ : MX2C
      port map(A => \data_temp[122]_net_1\, B => 
        \data_selected[154]\, S => \state[4]_net_1\, Y => N_723);
    
    \data_temp_RNO_2[95]\ : MX2C
      port map(A => data_f2_out(127), B => data_f3_out(127), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1720);
    
    \data_temp_RNO_0[100]\ : MX2C
      port map(A => \data_temp[100]_net_1\, B => 
        \data_selected[132]\, S => \state[4]_net_1\, Y => N_701);
    
    \data_temp_RNO[13]\ : NOR2A
      port map(A => \data_temp[45]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[13]\);
    
    \data_valid_and_ready[0]\ : OR2A
      port map(A => valid_out_0, B => ready_i_0(0), Y => 
        \data_valid_and_ready[0]_net_1\);
    
    \data_temp_RNO_3[97]\ : MX2C
      port map(A => data_f0_out(129), B => data_f1_out(129), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_785);
    
    \data[19]\ : DFN1C0
      port map(D => \data_5[19]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(19));
    
    \data_temp_RNO_0[84]\ : MX2C
      port map(A => \data_temp[116]_net_1\, B => 
        \data_selected[116]\, S => \state[4]_net_1\, Y => N_685);
    
    \time_wen[2]\ : DFN1E0P0
      port map(D => N_859, CLK => HCLK_c, PRE => HRESETn_c, E => 
        N_928, Q => time_wen(2));
    
    \data_temp[118]\ : DFN1C0
      port map(D => \data_temp_5[118]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[118]_net_1\);
    
    \data_temp_RNO[109]\ : NOR2A
      port map(A => N_863, B => N_710, Y => \data_temp_5[109]\);
    
    \data_temp_RNO_2[94]\ : MX2C
      port map(A => data_f2_out(126), B => data_f3_out(126), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1719);
    
    \data_temp_RNO_1[79]\ : MX2C
      port map(A => N_1732, B => N_809, S => N_1580_2, Y => 
        \data_selected[111]\);
    
    \data_temp_RNO_1[71]\ : MX2C
      port map(A => N_740, B => N_815, S => N_1580_3, Y => 
        \data_selected[103]\);
    
    \data_temp[105]\ : DFN1C0
      port map(D => \data_temp_5[105]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[105]_net_1\);
    
    \data_temp[42]\ : DFN1C0
      port map(D => N_237, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[42]_net_1\);
    
    \data_temp_RNO_0[65]\ : MX2C
      port map(A => \data_temp[97]_net_1\, B => 
        \data_selected[97]\, S => \state[4]_net_1\, Y => N_666);
    
    \data_temp_RNO[103]\ : NOR2A
      port map(A => N_863_2, B => N_704, Y => \data_temp_5[103]\);
    
    \data_temp_RNO_3[102]\ : MX2C
      port map(A => data_f0_out(134), B => data_f1_out(134), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_790);
    
    \data_temp_RNO_0[114]\ : MX2C
      port map(A => \data_temp[114]_net_1\, B => 
        \data_selected[146]\, S => \state[4]_net_1\, Y => N_715);
    
    \data[15]\ : DFN1C0
      port map(D => \data_5[15]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(15));
    
    \data_temp_RNO_0[111]\ : MX2C
      port map(A => \data_temp[111]_net_1\, B => 
        \data_selected[143]\, S => \state[4]_net_1\, Y => N_712);
    
    \data_RNO[26]\ : NOR2A
      port map(A => \data_temp[26]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[26]\);
    
    \data_temp[1]\ : DFN1C0
      port map(D => \data_temp_5[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[1]_net_1\);
    
    \data_temp_RNO_1[66]\ : MX2C
      port map(A => N_735, B => N_824, S => N_1580, Y => 
        \data_selected[98]\);
    
    \data_temp_RNO_1[89]\ : MX2C
      port map(A => N_1728, B => N_805, S => N_1580, Y => 
        \data_selected[121]\);
    
    \data_temp_RNO_1[81]\ : MX2C
      port map(A => N_1734, B => N_811, S => N_1580_2, Y => 
        \data_selected[113]\);
    
    \data_temp_RNO_0[64]\ : MX2C
      port map(A => \data_temp[96]_net_1\, B => 
        \data_selected[96]\, S => \state[4]_net_1\, Y => N_665);
    
    \data_temp_RNO_0[96]\ : MX2C
      port map(A => \data_temp[96]_net_1\, B => 
        \data_selected[128]\, S => \state[4]_net_1\, Y => N_697);
    
    \data_temp_RNO_1[58]\ : MX2C
      port map(A => N_741, B => N_830, S => N_1580_2, Y => 
        \data_selected[90]\);
    
    \data_temp_RNO_1[99]\ : MX2C
      port map(A => N_1724, B => N_787, S => N_1580, Y => 
        \data_selected[131]\);
    
    \data_temp_RNO_1[91]\ : MX2
      port map(A => data_f0_out(123), B => data_f1_out(123), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_793);
    
    \data_temp_RNO_1[63]\ : MX2C
      port map(A => N_746, B => N_821, S => N_1580_2, Y => 
        \data_selected[95]\);
    
    \data_temp_RNO_3[106]\ : MX2C
      port map(A => data_f0_out(138), B => data_f1_out(138), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_780);
    
    \data_temp_RNO[28]\ : NOR2A
      port map(A => \data_temp[60]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[28]\);
    
    \data_temp_RNO_1[32]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1685, 
        Y => N_865);
    
    \data_temp[41]\ : DFN1C0
      port map(D => N_235, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[41]_net_1\);
    
    \data_temp_RNO_2[78]\ : MX2C
      port map(A => data_f2_out(110), B => data_f3_out(110), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_733);
    
    \data_temp_RNO_0[93]\ : AO1D
      port map(A => N_912_i, B => N_795, C => N_902, Y => 
        \data_temp_5_i_0[93]\);
    
    \data_temp_RNO_0[50]\ : MX2C
      port map(A => \data_temp[82]_net_1\, B => 
        \data_selected[82]\, S => \state[4]_net_1\, Y => N_651);
    
    \data_temp_RNO[97]\ : NOR2A
      port map(A => N_863, B => N_698, Y => \data_temp_5[97]\);
    
    \data_temp_RNO_0[47]\ : MX2C
      port map(A => \data_temp[79]_net_1\, B => 
        \data_selected[79]\, S => \state[4]_net_1\, Y => N_648);
    
    \data_RNO[14]\ : NOR2A
      port map(A => \data_temp[14]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[14]\);
    
    \data_temp_RNO_3[40]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[72]_net_1\, 
        Y => N_1662);
    
    \data_temp[23]\ : DFN1C0
      port map(D => \data_temp_5[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[23]_net_1\);
    
    \data_temp_RNO_3[121]\ : MX2C
      port map(A => data_f0_out(153), B => data_f1_out(153), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1678);
    
    \data_temp_RNO_2[37]\ : MX2
      port map(A => data_f0_out(69), B => data_f1_out(69), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_851);
    
    \data_temp[19]\ : DFN1C0
      port map(D => \data_temp_5[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[19]_net_1\);
    
    \data_temp_RNO_2[48]\ : MX2C
      port map(A => data_f2_out(80), B => data_f3_out(80), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_759);
    
    \data_temp_RNO_1[75]\ : MX2C
      port map(A => N_730, B => N_819, S => N_1580_2, Y => 
        \data_selected[107]\);
    
    \data_valid_and_ready_0[0]\ : OR2A
      port map(A => valid_out_0, B => ready_i_0(0), Y => 
        \data_valid_and_ready_0[0]_net_1\);
    
    \data_temp_RNO[23]\ : NOR2A
      port map(A => \data_temp[55]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[23]\);
    
    \data_RNO[10]\ : NOR2A
      port map(A => \data_temp[10]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[10]\);
    
    \data_temp[60]\ : DFN1C0
      port map(D => \data_temp_5[60]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[60]_net_1\);
    
    \data_temp[53]\ : DFN1C0
      port map(D => \data_temp_5[53]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[53]_net_1\);
    
    \data_valid_and_ready_3[2]\ : OR2A
      port map(A => valid_out_2, B => ready_i_0(2), Y => 
        \data_valid_and_ready_3[2]_net_1\);
    
    \data_temp_RNO_3[76]\ : MX2C
      port map(A => data_f0_out(108), B => data_f1_out(108), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_806);
    
    \data_temp_RNO_1[74]\ : MX2C
      port map(A => N_729, B => N_818, S => N_1580_2, Y => 
        \data_selected[106]\);
    
    \data_temp_RNO_1[85]\ : MX2C
      port map(A => N_1738, B => N_801, S => N_1580_3, Y => 
        \data_selected[117]\);
    
    \data_wen_RNO[3]\ : OR2
      port map(A => \time_en_temp[3]_net_1\, B => 
        \state[4]_net_1\, Y => \data_wen_3[3]\);
    
    \data_temp_RNO_1[103]\ : MX2C
      port map(A => N_1714, B => N_791, S => N_1580_3, Y => 
        \data_selected[135]\);
    
    \data_RNO[8]\ : NOR2A
      port map(A => \data_temp[8]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[8]\);
    
    \data_temp_RNO_0[113]\ : MX2C
      port map(A => \data_temp[113]_net_1\, B => 
        \data_selected[145]\, S => \state[4]_net_1\, Y => N_714);
    
    \data_temp_RNO_0[76]\ : MX2C
      port map(A => \data_temp[108]_net_1\, B => 
        \data_selected[108]\, S => \state[4]_net_1\, Y => N_677);
    
    \data_temp_RNO[69]\ : NOR2A
      port map(A => N_863, B => N_670, Y => \data_temp_5[69]\);
    
    \data_temp_RNO_2[102]\ : MX2C
      port map(A => data_f2_out(134), B => data_f3_out(134), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1713);
    
    \data_temp_RNO_0[52]\ : MX2C
      port map(A => \data_temp[84]_net_1\, B => 
        \data_selected[84]\, S => \state[4]_net_1\, Y => N_653);
    
    \data_temp_RNO_1[125]\ : MX2
      port map(A => data_f0_out(157), B => data_f1_out(157), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1682);
    
    \data_RNO[9]\ : NOR2A
      port map(A => \data_temp[9]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[9]\);
    
    \data_temp_RNO_2[105]\ : MX2C
      port map(A => data_f2_out(137), B => data_f3_out(137), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1716);
    
    \data_temp_RNO_3[42]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[74]_net_1\, 
        Y => N_1668);
    
    \data_temp_RNO_1[111]\ : MX2C
      port map(A => N_1708, B => N_771, S => N_1580_2, Y => 
        \data_selected[143]\);
    
    \data_valid_ack[1]\ : DFN1E0C0
      port map(D => N_857, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_929, Q => valid_ack(1));
    
    \data_temp_RNO_3[73]\ : MX2C
      port map(A => data_f0_out(105), B => data_f1_out(105), S
         => \data_valid_and_ready_3[0]_net_1\, Y => N_817);
    
    \data_temp_RNO_1[84]\ : MX2C
      port map(A => N_1737, B => N_800, S => N_1580_3, Y => 
        \data_selected[116]\);
    
    \data_temp_RNO_1[95]\ : MX2C
      port map(A => N_1720, B => N_797, S => N_1580_1, Y => 
        \data_selected[127]\);
    
    \data_temp_RNO_1[40]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_765, 
        Y => N_1663);
    
    \data_temp[48]\ : DFN1C0
      port map(D => \data_temp_5[48]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[48]_net_1\);
    
    \data_temp_RNO[50]\ : NOR2A
      port map(A => N_863_1, B => N_651, Y => \data_temp_5[50]\);
    
    \data_temp[86]\ : DFN1C0
      port map(D => \data_temp_5[86]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[86]_net_1\);
    
    \state_RNI8220I_0[4]\ : NOR2A
      port map(A => \state[4]_net_1\, B => N_917, Y => N_857);
    
    \data_temp_RNO[3]\ : NOR2A
      port map(A => \data_temp[35]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[3]\);
    
    \data_temp_RNO_3[59]\ : MX2C
      port map(A => data_f0_out(91), B => data_f1_out(91), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_831);
    
    \data_temp_RNO_3[51]\ : MX2C
      port map(A => data_f0_out(83), B => data_f1_out(83), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_837);
    
    \data_temp_RNO[80]\ : NOR2A
      port map(A => N_863_1, B => N_681, Y => \data_temp_5[80]\);
    
    \data_temp_RNO_3[125]\ : MX2
      port map(A => data_f2_out(157), B => data_f3_out(157), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1694);
    
    \data_temp_RNO_3[69]\ : MX2C
      port map(A => data_f0_out(101), B => data_f1_out(101), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_813);
    
    \data_temp_RNO_3[61]\ : MX2C
      port map(A => data_f0_out(93), B => data_f1_out(93), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_833);
    
    \data_temp_RNO_0[73]\ : MX2C
      port map(A => \data_temp[105]_net_1\, B => 
        \data_selected[105]\, S => \state[4]_net_1\, Y => N_674);
    
    \data_RNO[15]\ : NOR2A
      port map(A => \data_temp[15]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[15]\);
    
    \data_temp_RNO_3[89]\ : MX2C
      port map(A => data_f0_out(121), B => data_f1_out(121), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_805);
    
    \data_temp_RNO_3[81]\ : MX2C
      port map(A => data_f0_out(113), B => data_f1_out(113), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_811);
    
    \data_temp_RNO[66]\ : NOR2A
      port map(A => N_863, B => N_667, Y => \data_temp_5[66]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \data_temp_RNO_3[109]\ : MX2C
      port map(A => data_f0_out(141), B => data_f1_out(141), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_783);
    
    \data_temp[116]\ : DFN1C0
      port map(D => \data_temp_5[116]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[116]_net_1\);
    
    \data_temp_RNO_1[94]\ : MX2C
      port map(A => N_1719, B => N_796, S => N_1580_1, Y => 
        \data_selected[126]\);
    
    \data_temp_RNO[11]\ : NOR2A
      port map(A => \data_temp[43]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[11]\);
    
    \data_temp_RNO_1[126]\ : MX2C
      port map(A => N_1695, B => N_1683, S => N_1580_1, Y => 
        \data_selected[158]\);
    
    \data_temp_RNO_4[36]\ : MX2
      port map(A => data_f2_out(68), B => data_f3_out(68), S => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_1689);
    
    \data_RNO[29]\ : NOR2A
      port map(A => \data_temp[29]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[29]\);
    
    \state[3]\ : DFN1C0
      port map(D => state_0_sqmuxa_i_i, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \state[3]_net_1\);
    
    \data_temp_RNO[12]\ : NOR2A
      port map(A => \data_temp[44]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[12]\);
    
    \data_temp[47]\ : DFN1C0
      port map(D => \data_temp_5[47]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[47]_net_1\);
    
    \data_valid_ack_RNO[2]\ : INV
      port map(A => N_859, Y => N_859_i);
    
    \data_RNO[30]\ : NOR2A
      port map(A => \data_temp[30]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[30]\);
    
    \data_temp_RNO_4[33]\ : MX2
      port map(A => data_f2_out(65), B => data_f3_out(65), S => 
        \data_valid_and_ready_0[2]_net_1\, Y => N_1686);
    
    \data_temp_RNO_3[90]\ : MX2C
      port map(A => data_f0_out(122), B => data_f1_out(122), S
         => \data_valid_and_ready_1[0]_net_1\, Y => N_792);
    
    \data_temp_RNO_1[42]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_767, 
        Y => N_1669);
    
    \data_temp_RNO_2[121]\ : MX2C
      port map(A => data_f2_out(153), B => data_f3_out(153), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1690);
    
    \data_temp[33]\ : DFN1C0
      port map(D => N_219, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \data_temp[33]_net_1\);
    
    \data_temp[20]\ : DFN1C0
      port map(D => \data_temp_5[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[20]_net_1\);
    
    \data_temp_RNO_2[106]\ : MX2C
      port map(A => data_f2_out(138), B => data_f3_out(138), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1717);
    
    \data_temp_RNIERBC[125]\ : OR2
      port map(A => \state[4]_net_1\, B => \data_temp[125]_net_1\, 
        Y => N_914);
    
    \data[24]\ : DFN1C0
      port map(D => \data_5[24]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(24));
    
    \data_temp_RNO[95]\ : NOR2A
      port map(A => N_863_0, B => N_696, Y => \data_temp_5[95]\);
    
    \data_temp_RNO[14]\ : NOR2A
      port map(A => \data_temp[46]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[14]\);
    
    \data_temp_RNO_2[89]\ : MX2C
      port map(A => data_f2_out(121), B => data_f3_out(121), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1728);
    
    \data_temp_RNO_2[81]\ : MX2C
      port map(A => data_f2_out(113), B => data_f3_out(113), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1734);
    
    \data_temp_RNO_3[39]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[71]_net_1\, 
        Y => N_1659);
    
    \data_temp[50]\ : DFN1C0
      port map(D => \data_temp_5[50]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[50]_net_1\);
    
    \data_temp_RNO_3[55]\ : MX2C
      port map(A => data_f0_out(87), B => data_f1_out(87), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_827);
    
    \data_temp_RNO_0[86]\ : MX2C
      port map(A => \data_temp[118]_net_1\, B => 
        \data_selected[118]\, S => \state[4]_net_1\, Y => N_687);
    
    \data[1]\ : DFN1C0
      port map(D => \data_5[1]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(1));
    
    \data_valid_and_ready_2[2]\ : OR2A
      port map(A => valid_out_2, B => ready_i_0(2), Y => 
        \data_valid_and_ready_2[2]_net_1\);
    
    \data_temp_RNO_3[65]\ : MX2C
      port map(A => data_f0_out(97), B => data_f1_out(97), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_823);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \data_valid_and_ready[1]\ : NOR2
      port map(A => valid_out_i(1), B => ready_i_0(1), Y => 
        \data_valid_and_ready[1]_net_1\);
    
    \data_temp_RNO_3[85]\ : MX2C
      port map(A => data_f0_out(117), B => data_f1_out(117), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_801);
    
    \state_RNO[4]\ : OA1B
      port map(A => N_1306, B => \state[0]_net_1\, C => 
        \state_ns_i_i_a2_1[0]\, Y => N_861);
    
    \data_temp_RNO_2[96]\ : MX2C
      port map(A => data_f2_out(128), B => data_f3_out(128), S
         => \data_valid_and_ready_1[2]_net_1\, Y => N_1721);
    
    \data[9]\ : DFN1C0
      port map(D => \data_5[9]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(9));
    
    \data_temp_RNO_3[123]\ : MX2
      port map(A => data_f2_out(155), B => data_f3_out(155), S
         => \data_valid_and_ready_0[2]_net_1\, Y => N_1692);
    
    \data_valid_and_ready[2]\ : OR2A
      port map(A => valid_out_2, B => ready_i_0(2), Y => 
        \data_valid_and_ready[2]_net_1\);
    
    \data_temp_RNO_3[54]\ : MX2C
      port map(A => data_f0_out(86), B => data_f1_out(86), S => 
        \data_valid_and_ready[0]_net_1\, Y => N_840);
    
    \data_temp_RNO_1[124]\ : MX2
      port map(A => data_f0_out(156), B => data_f1_out(156), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1681);
    
    \data_temp_RNO_3[92]\ : MX2
      port map(A => data_f2_out(124), B => data_f3_out(124), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1731);
    
    \data_temp_RNO_3[64]\ : MX2C
      port map(A => data_f0_out(96), B => data_f1_out(96), S => 
        \data_valid_and_ready_3[0]_net_1\, Y => N_822);
    
    \data_temp_RNO_1[57]\ : MX2C
      port map(A => N_754, B => N_829, S => N_1580_1, Y => 
        \data_selected[89]\);
    
    \data_temp_RNO_2[69]\ : MX2C
      port map(A => data_f2_out(101), B => data_f3_out(101), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_738);
    
    \data_temp_RNO_2[61]\ : MX2C
      port map(A => data_f2_out(93), B => data_f3_out(93), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_744);
    
    \data[17]\ : DFN1C0
      port map(D => \data_5[17]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(17));
    
    \data_temp_RNO_3[84]\ : MX2C
      port map(A => data_f0_out(116), B => data_f1_out(116), S
         => \data_valid_and_ready_2[0]_net_1\, Y => N_800);
    
    \data_temp_RNO_0[83]\ : MX2C
      port map(A => \data_temp[115]_net_1\, B => 
        \data_selected[115]\, S => \state[4]_net_1\, Y => N_684);
    
    \data_temp_RNO_2[58]\ : MX2C
      port map(A => data_f2_out(90), B => data_f3_out(90), S => 
        \data_valid_and_ready_3[2]_net_1\, Y => N_741);
    
    \data[20]\ : DFN1C0
      port map(D => \data_5[20]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => wdata(20));
    
    \data_temp_RNO_2[93]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_0, C => N_1718, 
        Y => N_902);
    
    \data_RNO[6]\ : NOR2A
      port map(A => \data_temp[6]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[6]\);
    
    \data_RNO[3]\ : NOR2A
      port map(A => \data_temp[3]_net_1\, B => \state[4]_net_1\, 
        Y => \data_5[3]\);
    
    \data_temp_RNO_2[77]\ : MX2C
      port map(A => data_f2_out(109), B => data_f3_out(109), S
         => \data_valid_and_ready_3[2]_net_1\, Y => N_732);
    
    \data_temp_RNO_0[66]\ : MX2C
      port map(A => \data_temp[98]_net_1\, B => 
        \data_selected[98]\, S => \state[4]_net_1\, Y => N_667);
    
    \data_temp_RNO[21]\ : NOR2A
      port map(A => \data_temp[53]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[21]\);
    
    \data_wen[0]\ : DFN1E0P0
      port map(D => \data_wen_3[0]\, CLK => HCLK_c, PRE => 
        HRESETn_c, E => N_928, Q => data_wen(0));
    
    \data_temp_RNO_0[104]\ : MX2C
      port map(A => \data_temp[104]_net_1\, B => 
        \data_selected[136]\, S => \state[4]_net_1\, Y => N_705);
    
    \data_temp_RNO_4[40]\ : MX2
      port map(A => data_f2_out(72), B => data_f3_out(72), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_765);
    
    \data_temp_RNO_2[47]\ : MX2C
      port map(A => data_f2_out(79), B => data_f3_out(79), S => 
        \data_valid_and_ready[2]_net_1\, Y => N_758);
    
    \data_temp_RNO_0[101]\ : MX2C
      port map(A => \data_temp[101]_net_1\, B => 
        \data_selected[133]\, S => \state[4]_net_1\, Y => N_702);
    
    \data_temp_RNO_0[40]\ : AO1D
      port map(A => N_912_i, B => N_854, C => N_1662, Y => 
        \data_temp_5_i_0[40]\);
    
    \data_temp_RNO_0[38]\ : AO1D
      port map(A => N_912_i, B => N_852, C => N_1656, Y => 
        \data_temp_5_i_0[38]\);
    
    \state_RNIIO749[4]\ : OR2A
      port map(A => \state[4]_net_1\, B => 
        \data_valid_and_ready_0[0]_net_1\, Y => \time_wen_3[0]\);
    
    \data_temp_RNO[67]\ : NOR2A
      port map(A => N_863, B => N_668, Y => \data_temp_5[67]\);
    
    \data_temp_RNO[22]\ : NOR2A
      port map(A => \data_temp[54]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[22]\);
    
    \data_temp_RNO[79]\ : NOR2A
      port map(A => N_863_2, B => N_680, Y => \data_temp_5[79]\);
    
    \data_temp[66]\ : DFN1C0
      port map(D => \data_temp_5[66]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[66]_net_1\);
    
    \data_temp_RNO_2[85]\ : MX2C
      port map(A => data_f2_out(117), B => data_f3_out(117), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1738);
    
    \data_temp_RNO_2[123]\ : NOR3A
      port map(A => \state[4]_net_1\, B => N_1580_1, C => N_1692, 
        Y => N_910);
    
    \data_temp_RNO_0[63]\ : MX2C
      port map(A => \data_temp[95]_net_1\, B => 
        \data_selected[95]\, S => \state[4]_net_1\, Y => N_664);
    
    \data_temp_RNO_3[35]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[67]_net_1\, 
        Y => N_873);
    
    \data_temp[84]\ : DFN1C0
      port map(D => \data_temp_5[84]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[84]_net_1\);
    
    \data_temp[45]\ : DFN1C0
      port map(D => \data_temp_5[45]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[45]_net_1\);
    
    \data_valid_ack[2]\ : DFN1E0C0
      port map(D => N_859_i, CLK => HCLK_c, CLR => HRESETn_c, E
         => N_929, Q => valid_ack(2));
    
    \data_temp[73]\ : DFN1C0
      port map(D => \data_temp_5[73]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[73]_net_1\);
    
    \data_temp_RNO_3[118]\ : MX2C
      port map(A => data_f0_out(150), B => data_f1_out(150), S
         => \data_valid_and_ready_0[0]_net_1\, Y => N_1675);
    
    \data_temp_RNO_2[84]\ : MX2C
      port map(A => data_f2_out(116), B => data_f3_out(116), S
         => \data_valid_and_ready_2[2]_net_1\, Y => N_1737);
    
    \data_temp_RNO[76]\ : NOR2A
      port map(A => N_863_1, B => N_677, Y => \data_temp_5[76]\);
    
    \data_temp_RNO_3[34]\ : NOR2
      port map(A => \state[4]_net_1\, B => \data_temp[66]_net_1\, 
        Y => N_870);
    
    \data_temp[113]\ : DFN1C0
      port map(D => \data_temp_5[113]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[113]_net_1\);
    
    \data_temp_RNO[24]\ : NOR2A
      port map(A => \data_temp[56]_net_1\, B => \state[4]_net_1\, 
        Y => \data_temp_5[24]\);
    
    \data_temp[30]\ : DFN1C0
      port map(D => \data_temp_5[30]\, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => \data_temp[30]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_waveform is

    port( status_full_ack    : in    std_logic_vector(3 downto 0);
          hburst_c           : out   std_logic_vector(2 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          hsize_c            : out   std_logic_vector(1 downto 0);
          AHB_Master_In_c_5  : in    std_logic;
          AHB_Master_In_c_4  : in    std_logic;
          AHB_Master_In_c_0  : in    std_logic;
          AHB_Master_In_c_3  : in    std_logic;
          haddr_c            : out   std_logic_vector(31 downto 0);
          nb_burst_available : in    std_logic_vector(10 downto 0);
          status_full_err    : out   std_logic_vector(3 downto 0);
          status_full        : out   std_logic_vector(3 downto 0);
          addr_data_f3       : in    std_logic_vector(31 downto 0);
          addr_data_f2       : in    std_logic_vector(31 downto 0);
          addr_data_f1       : in    std_logic_vector(31 downto 0);
          addr_data_f0       : in    std_logic_vector(31 downto 0);
          hwdata_c           : out   std_logic_vector(31 downto 0);
          status_new_err     : out   std_logic_vector(3 downto 0);
          sample_f3_wdata    : in    std_logic_vector(95 downto 0);
          sample_f2_wdata    : in    std_logic_vector(95 downto 0);
          sample_f1_15       : in    std_logic;
          sample_f1_47       : in    std_logic;
          sample_f1_14       : in    std_logic;
          sample_f1_46       : in    std_logic;
          sample_f1_13       : in    std_logic;
          sample_f1_45       : in    std_logic;
          sample_f1_12       : in    std_logic;
          sample_f1_44       : in    std_logic;
          sample_f1_60       : in    std_logic;
          sample_f1_59       : in    std_logic;
          sample_f1_58       : in    std_logic;
          sample_f1_57       : in    std_logic;
          sample_f1_56       : in    std_logic;
          sample_f1_55       : in    std_logic;
          sample_f1_54       : in    std_logic;
          sample_f1_53       : in    std_logic;
          sample_f1_52       : in    std_logic;
          sample_f1_51       : in    std_logic;
          sample_f1_50       : in    std_logic;
          sample_f1_49       : in    std_logic;
          sample_f1_48       : in    std_logic;
          sample_f1_4        : in    std_logic;
          sample_f1_36       : in    std_logic;
          sample_f1_3        : in    std_logic;
          sample_f1_35       : in    std_logic;
          sample_f1_2        : in    std_logic;
          sample_f1_34       : in    std_logic;
          sample_f1_1        : in    std_logic;
          sample_f1_33       : in    std_logic;
          sample_f1_0        : in    std_logic;
          sample_f1_32       : in    std_logic;
          sample_f1_63       : in    std_logic;
          sample_f1_62       : in    std_logic;
          sample_f1_61       : in    std_logic;
          sample_f1_11       : in    std_logic;
          sample_f1_43       : in    std_logic;
          sample_f1_10       : in    std_logic;
          sample_f1_42       : in    std_logic;
          sample_f1_9        : in    std_logic;
          sample_f1_41       : in    std_logic;
          sample_f1_8        : in    std_logic;
          sample_f1_40       : in    std_logic;
          sample_f1_7        : in    std_logic;
          sample_f1_39       : in    std_logic;
          sample_f1_6        : in    std_logic;
          sample_f1_38       : in    std_logic;
          sample_f1_5        : in    std_logic;
          sample_f1_37       : in    std_logic;
          sample_f1_wdata_0  : in    std_logic;
          sample_f1_wdata_1  : in    std_logic;
          sample_f1_wdata_2  : in    std_logic;
          sample_f1_wdata_3  : in    std_logic;
          sample_f1_wdata_4  : in    std_logic;
          sample_f1_wdata_5  : in    std_logic;
          sample_f1_wdata_6  : in    std_logic;
          sample_f1_wdata_7  : in    std_logic;
          sample_f1_wdata_8  : in    std_logic;
          sample_f1_wdata_9  : in    std_logic;
          sample_f1_wdata_10 : in    std_logic;
          sample_f1_wdata_11 : in    std_logic;
          sample_f1_wdata_12 : in    std_logic;
          sample_f1_wdata_13 : in    std_logic;
          sample_f1_wdata_14 : in    std_logic;
          sample_f1_wdata_15 : in    std_logic;
          sample_f1_wdata_48 : in    std_logic;
          sample_f1_wdata_49 : in    std_logic;
          sample_f1_wdata_50 : in    std_logic;
          sample_f1_wdata_51 : in    std_logic;
          sample_f1_wdata_52 : in    std_logic;
          sample_f1_wdata_53 : in    std_logic;
          sample_f1_wdata_54 : in    std_logic;
          sample_f1_wdata_55 : in    std_logic;
          sample_f1_wdata_56 : in    std_logic;
          sample_f1_wdata_57 : in    std_logic;
          sample_f1_wdata_58 : in    std_logic;
          sample_f1_wdata_59 : in    std_logic;
          sample_f1_wdata_60 : in    std_logic;
          sample_f1_wdata_61 : in    std_logic;
          sample_f1_wdata_62 : in    std_logic;
          sample_f1_wdata_63 : in    std_logic;
          sample_f1_wdata_64 : in    std_logic;
          sample_f1_wdata_65 : in    std_logic;
          sample_f1_wdata_66 : in    std_logic;
          sample_f1_wdata_67 : in    std_logic;
          sample_f1_wdata_68 : in    std_logic;
          sample_f1_wdata_69 : in    std_logic;
          sample_f1_wdata_70 : in    std_logic;
          sample_f1_wdata_71 : in    std_logic;
          sample_f1_wdata_72 : in    std_logic;
          sample_f1_wdata_73 : in    std_logic;
          sample_f1_wdata_74 : in    std_logic;
          sample_f1_wdata_75 : in    std_logic;
          sample_f1_wdata_76 : in    std_logic;
          sample_f1_wdata_77 : in    std_logic;
          sample_f1_wdata_78 : in    std_logic;
          sample_f1_wdata_79 : in    std_logic;
          sample_f1_wdata_80 : in    std_logic;
          sample_f1_wdata_81 : in    std_logic;
          sample_f1_wdata_82 : in    std_logic;
          sample_f1_wdata_83 : in    std_logic;
          sample_f1_wdata_84 : in    std_logic;
          sample_f1_wdata_85 : in    std_logic;
          sample_f1_wdata_86 : in    std_logic;
          sample_f1_wdata_87 : in    std_logic;
          sample_f1_wdata_88 : in    std_logic;
          sample_f1_wdata_89 : in    std_logic;
          sample_f1_wdata_90 : in    std_logic;
          sample_f1_wdata_91 : in    std_logic;
          sample_f1_wdata_92 : in    std_logic;
          sample_f1_wdata_93 : in    std_logic;
          sample_f1_wdata_94 : in    std_logic;
          sample_f1_wdata_95 : in    std_logic;
          sample_f0_15       : in    std_logic;
          sample_f0_47       : in    std_logic;
          sample_f0_14       : in    std_logic;
          sample_f0_46       : in    std_logic;
          sample_f0_13       : in    std_logic;
          sample_f0_45       : in    std_logic;
          sample_f0_12       : in    std_logic;
          sample_f0_44       : in    std_logic;
          sample_f0_60       : in    std_logic;
          sample_f0_59       : in    std_logic;
          sample_f0_58       : in    std_logic;
          sample_f0_57       : in    std_logic;
          sample_f0_56       : in    std_logic;
          sample_f0_55       : in    std_logic;
          sample_f0_54       : in    std_logic;
          sample_f0_53       : in    std_logic;
          sample_f0_52       : in    std_logic;
          sample_f0_51       : in    std_logic;
          sample_f0_50       : in    std_logic;
          sample_f0_49       : in    std_logic;
          sample_f0_48       : in    std_logic;
          sample_f0_4        : in    std_logic;
          sample_f0_36       : in    std_logic;
          sample_f0_3        : in    std_logic;
          sample_f0_35       : in    std_logic;
          sample_f0_2        : in    std_logic;
          sample_f0_34       : in    std_logic;
          sample_f0_1        : in    std_logic;
          sample_f0_33       : in    std_logic;
          sample_f0_0        : in    std_logic;
          sample_f0_32       : in    std_logic;
          sample_f0_63       : in    std_logic;
          sample_f0_62       : in    std_logic;
          sample_f0_61       : in    std_logic;
          sample_f0_11       : in    std_logic;
          sample_f0_43       : in    std_logic;
          sample_f0_10       : in    std_logic;
          sample_f0_42       : in    std_logic;
          sample_f0_9        : in    std_logic;
          sample_f0_41       : in    std_logic;
          sample_f0_8        : in    std_logic;
          sample_f0_40       : in    std_logic;
          sample_f0_7        : in    std_logic;
          sample_f0_39       : in    std_logic;
          sample_f0_6        : in    std_logic;
          sample_f0_38       : in    std_logic;
          sample_f0_5        : in    std_logic;
          sample_f0_37       : in    std_logic;
          sample_f0_wdata_0  : in    std_logic;
          sample_f0_wdata_1  : in    std_logic;
          sample_f0_wdata_2  : in    std_logic;
          sample_f0_wdata_3  : in    std_logic;
          sample_f0_wdata_4  : in    std_logic;
          sample_f0_wdata_5  : in    std_logic;
          sample_f0_wdata_6  : in    std_logic;
          sample_f0_wdata_7  : in    std_logic;
          sample_f0_wdata_8  : in    std_logic;
          sample_f0_wdata_9  : in    std_logic;
          sample_f0_wdata_10 : in    std_logic;
          sample_f0_wdata_11 : in    std_logic;
          sample_f0_wdata_12 : in    std_logic;
          sample_f0_wdata_13 : in    std_logic;
          sample_f0_wdata_14 : in    std_logic;
          sample_f0_wdata_15 : in    std_logic;
          sample_f0_wdata_48 : in    std_logic;
          sample_f0_wdata_49 : in    std_logic;
          sample_f0_wdata_50 : in    std_logic;
          sample_f0_wdata_51 : in    std_logic;
          sample_f0_wdata_52 : in    std_logic;
          sample_f0_wdata_53 : in    std_logic;
          sample_f0_wdata_54 : in    std_logic;
          sample_f0_wdata_55 : in    std_logic;
          sample_f0_wdata_56 : in    std_logic;
          sample_f0_wdata_57 : in    std_logic;
          sample_f0_wdata_58 : in    std_logic;
          sample_f0_wdata_59 : in    std_logic;
          sample_f0_wdata_60 : in    std_logic;
          sample_f0_wdata_61 : in    std_logic;
          sample_f0_wdata_62 : in    std_logic;
          sample_f0_wdata_63 : in    std_logic;
          sample_f0_wdata_64 : in    std_logic;
          sample_f0_wdata_65 : in    std_logic;
          sample_f0_wdata_66 : in    std_logic;
          sample_f0_wdata_67 : in    std_logic;
          sample_f0_wdata_68 : in    std_logic;
          sample_f0_wdata_69 : in    std_logic;
          sample_f0_wdata_70 : in    std_logic;
          sample_f0_wdata_71 : in    std_logic;
          sample_f0_wdata_72 : in    std_logic;
          sample_f0_wdata_73 : in    std_logic;
          sample_f0_wdata_74 : in    std_logic;
          sample_f0_wdata_75 : in    std_logic;
          sample_f0_wdata_76 : in    std_logic;
          sample_f0_wdata_77 : in    std_logic;
          sample_f0_wdata_78 : in    std_logic;
          sample_f0_wdata_79 : in    std_logic;
          sample_f0_wdata_80 : in    std_logic;
          sample_f0_wdata_81 : in    std_logic;
          sample_f0_wdata_82 : in    std_logic;
          sample_f0_wdata_83 : in    std_logic;
          sample_f0_wdata_84 : in    std_logic;
          sample_f0_wdata_85 : in    std_logic;
          sample_f0_wdata_86 : in    std_logic;
          sample_f0_wdata_87 : in    std_logic;
          sample_f0_wdata_88 : in    std_logic;
          sample_f0_wdata_89 : in    std_logic;
          sample_f0_wdata_90 : in    std_logic;
          sample_f0_wdata_91 : in    std_logic;
          sample_f0_wdata_92 : in    std_logic;
          sample_f0_wdata_93 : in    std_logic;
          sample_f0_wdata_94 : in    std_logic;
          sample_f0_wdata_95 : in    std_logic;
          delta_f2_f1        : in    std_logic_vector(9 downto 0);
          delta_snapshot     : in    std_logic_vector(15 downto 0);
          delta_f2_f0        : in    std_logic_vector(9 downto 0);
          nb_snapshot_param  : in    std_logic_vector(10 downto 0);
          hwrite_c           : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          N_43               : out   std_logic;
          lpp_waveform_GND   : in    std_logic;
          lpp_waveform_VCC   : in    std_logic;
          sample_f3_val      : in    std_logic;
          enable_f3          : in    std_logic;
          burst_f2           : in    std_logic;
          enable_f2          : in    std_logic;
          sample_f1_val_0    : in    std_logic;
          burst_f1           : in    std_logic;
          enable_f1          : in    std_logic;
          data_shaping_R1_0  : in    std_logic;
          data_shaping_R1    : in    std_logic;
          burst_f0           : in    std_logic;
          data_shaping_R0_0  : in    std_logic;
          data_shaping_R0    : in    std_logic;
          enable_f0          : in    std_logic;
          coarse_time_0_c    : in    std_logic;
          sample_f2_val      : in    std_logic;
          sample_f0_val_0    : in    std_logic;
          HCLK_c             : in    std_logic;
          HRESETn_c          : in    std_logic
        );

end lpp_waveform;

architecture DEF_ARCH of lpp_waveform is 

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1
    port( sample_f1_wdata_95 : in    std_logic := 'U';
          sample_f1_wdata_94 : in    std_logic := 'U';
          sample_f1_wdata_93 : in    std_logic := 'U';
          sample_f1_wdata_92 : in    std_logic := 'U';
          sample_f1_wdata_91 : in    std_logic := 'U';
          sample_f1_wdata_90 : in    std_logic := 'U';
          sample_f1_wdata_89 : in    std_logic := 'U';
          sample_f1_wdata_88 : in    std_logic := 'U';
          sample_f1_wdata_87 : in    std_logic := 'U';
          sample_f1_wdata_86 : in    std_logic := 'U';
          sample_f1_wdata_85 : in    std_logic := 'U';
          sample_f1_wdata_84 : in    std_logic := 'U';
          sample_f1_wdata_83 : in    std_logic := 'U';
          sample_f1_wdata_82 : in    std_logic := 'U';
          sample_f1_wdata_81 : in    std_logic := 'U';
          sample_f1_wdata_80 : in    std_logic := 'U';
          sample_f1_wdata_79 : in    std_logic := 'U';
          sample_f1_wdata_78 : in    std_logic := 'U';
          sample_f1_wdata_77 : in    std_logic := 'U';
          sample_f1_wdata_76 : in    std_logic := 'U';
          sample_f1_wdata_75 : in    std_logic := 'U';
          sample_f1_wdata_74 : in    std_logic := 'U';
          sample_f1_wdata_73 : in    std_logic := 'U';
          sample_f1_wdata_72 : in    std_logic := 'U';
          sample_f1_wdata_71 : in    std_logic := 'U';
          sample_f1_wdata_70 : in    std_logic := 'U';
          sample_f1_wdata_69 : in    std_logic := 'U';
          sample_f1_wdata_68 : in    std_logic := 'U';
          sample_f1_wdata_67 : in    std_logic := 'U';
          sample_f1_wdata_66 : in    std_logic := 'U';
          sample_f1_wdata_65 : in    std_logic := 'U';
          sample_f1_wdata_64 : in    std_logic := 'U';
          sample_f1_wdata_63 : in    std_logic := 'U';
          sample_f1_wdata_62 : in    std_logic := 'U';
          sample_f1_wdata_61 : in    std_logic := 'U';
          sample_f1_wdata_60 : in    std_logic := 'U';
          sample_f1_wdata_59 : in    std_logic := 'U';
          sample_f1_wdata_58 : in    std_logic := 'U';
          sample_f1_wdata_57 : in    std_logic := 'U';
          sample_f1_wdata_56 : in    std_logic := 'U';
          sample_f1_wdata_55 : in    std_logic := 'U';
          sample_f1_wdata_54 : in    std_logic := 'U';
          sample_f1_wdata_53 : in    std_logic := 'U';
          sample_f1_wdata_52 : in    std_logic := 'U';
          sample_f1_wdata_51 : in    std_logic := 'U';
          sample_f1_wdata_50 : in    std_logic := 'U';
          sample_f1_wdata_49 : in    std_logic := 'U';
          sample_f1_wdata_48 : in    std_logic := 'U';
          sample_f1_wdata_15 : in    std_logic := 'U';
          sample_f1_wdata_14 : in    std_logic := 'U';
          sample_f1_wdata_13 : in    std_logic := 'U';
          sample_f1_wdata_12 : in    std_logic := 'U';
          sample_f1_wdata_11 : in    std_logic := 'U';
          sample_f1_wdata_10 : in    std_logic := 'U';
          sample_f1_wdata_9  : in    std_logic := 'U';
          sample_f1_wdata_8  : in    std_logic := 'U';
          sample_f1_wdata_7  : in    std_logic := 'U';
          sample_f1_wdata_6  : in    std_logic := 'U';
          sample_f1_wdata_5  : in    std_logic := 'U';
          sample_f1_wdata_4  : in    std_logic := 'U';
          sample_f1_wdata_3  : in    std_logic := 'U';
          sample_f1_wdata_2  : in    std_logic := 'U';
          sample_f1_wdata_1  : in    std_logic := 'U';
          sample_f1_wdata_0  : in    std_logic := 'U';
          data_f1_out        : out   std_logic_vector(159 downto 64);
          nb_snapshot_param  : in    std_logic_vector(0 to 0) := (others => 'U');
          sample_f1_37       : in    std_logic := 'U';
          sample_f1_5        : in    std_logic := 'U';
          sample_f1_38       : in    std_logic := 'U';
          sample_f1_6        : in    std_logic := 'U';
          sample_f1_39       : in    std_logic := 'U';
          sample_f1_7        : in    std_logic := 'U';
          sample_f1_40       : in    std_logic := 'U';
          sample_f1_8        : in    std_logic := 'U';
          sample_f1_41       : in    std_logic := 'U';
          sample_f1_9        : in    std_logic := 'U';
          sample_f1_42       : in    std_logic := 'U';
          sample_f1_10       : in    std_logic := 'U';
          sample_f1_43       : in    std_logic := 'U';
          sample_f1_11       : in    std_logic := 'U';
          sample_f1_61       : in    std_logic := 'U';
          sample_f1_62       : in    std_logic := 'U';
          sample_f1_63       : in    std_logic := 'U';
          sample_f1_32       : in    std_logic := 'U';
          sample_f1_0        : in    std_logic := 'U';
          sample_f1_33       : in    std_logic := 'U';
          sample_f1_1        : in    std_logic := 'U';
          sample_f1_34       : in    std_logic := 'U';
          sample_f1_2        : in    std_logic := 'U';
          sample_f1_35       : in    std_logic := 'U';
          sample_f1_3        : in    std_logic := 'U';
          sample_f1_36       : in    std_logic := 'U';
          sample_f1_4        : in    std_logic := 'U';
          sample_f1_48       : in    std_logic := 'U';
          sample_f1_49       : in    std_logic := 'U';
          sample_f1_50       : in    std_logic := 'U';
          sample_f1_51       : in    std_logic := 'U';
          sample_f1_52       : in    std_logic := 'U';
          sample_f1_53       : in    std_logic := 'U';
          sample_f1_54       : in    std_logic := 'U';
          sample_f1_55       : in    std_logic := 'U';
          sample_f1_56       : in    std_logic := 'U';
          sample_f1_57       : in    std_logic := 'U';
          sample_f1_58       : in    std_logic := 'U';
          sample_f1_59       : in    std_logic := 'U';
          sample_f1_60       : in    std_logic := 'U';
          sample_f1_44       : in    std_logic := 'U';
          sample_f1_12       : in    std_logic := 'U';
          sample_f1_45       : in    std_logic := 'U';
          sample_f1_13       : in    std_logic := 'U';
          sample_f1_46       : in    std_logic := 'U';
          sample_f1_14       : in    std_logic := 'U';
          sample_f1_47       : in    std_logic := 'U';
          sample_f1_15       : in    std_logic := 'U';
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          data_f1_out_valid  : out   std_logic;
          N_4                : in    std_logic := 'U';
          I_38_4             : in    std_logic := 'U';
          I_24_4             : in    std_logic := 'U';
          I_20_12            : in    std_logic := 'U';
          I_13_20            : in    std_logic := 'U';
          I_45_4             : in    std_logic := 'U';
          I_9_20             : in    std_logic := 'U';
          I_5_20             : in    std_logic := 'U';
          I_52_4             : in    std_logic := 'U';
          data_shaping_R1    : in    std_logic := 'U';
          data_shaping_R1_0  : in    std_logic := 'U';
          I_56_4             : in    std_logic := 'U';
          I_31_5             : in    std_logic := 'U';
          enable_f1          : in    std_logic := 'U';
          burst_f1           : in    std_logic := 'U';
          sample_f1_val_0    : in    std_logic := 'U';
          start_snapshot_f1  : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_snapshot_controler
    port( delta_f2_f0       : in    std_logic_vector(9 downto 0) := (others => 'U');
          delta_snapshot    : in    std_logic_vector(15 downto 0) := (others => 'U');
          delta_f2_f1       : in    std_logic_vector(9 downto 0) := (others => 'U');
          start_snapshot_f2 : out   std_logic;
          start_snapshot_f1 : out   std_logic;
          start_snapshot_f0 : out   std_logic;
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          sample_f0_val_0   : in    std_logic := 'U';
          sample_f2_val     : in    std_logic := 'U';
          coarse_time_0_c   : in    std_logic := 'U'
        );
  end component;

  component 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\
    port( status_new_err    : out   std_logic_vector(3 to 3);
          valid_ack         : in    std_logic_vector(3 to 3) := (others => 'U');
          valid_out         : out   std_logic_vector(3 to 3);
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f3_out_valid : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\
    port( status_new_err    : out   std_logic_vector(1 to 1);
          valid_out_i       : out   std_logic_vector(1 to 1);
          valid_ack         : in    std_logic_vector(1 to 1) := (others => 'U');
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f1_out_valid : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component lpp_waveform_burst
    port( sample_f3_wdata   : in    std_logic_vector(95 downto 0) := (others => 'U');
          data_f3_out       : out   std_logic_vector(159 downto 64);
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f3_out_valid : out   std_logic;
          enable_f3         : in    std_logic := 'U';
          sample_f3_val     : in    std_logic := 'U'
        );
  end component;

  component 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\
    port( status_new_err    : out   std_logic_vector(2 to 2);
          valid_ack         : in    std_logic_vector(2 to 2) := (others => 'U');
          valid_out         : out   std_logic_vector(2 to 2);
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f2_out_valid : in    std_logic := 'U'
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\
    port( status_new_err    : out   std_logic_vector(0 to 0);
          valid_ack         : in    std_logic_vector(0 to 0) := (others => 'U');
          valid_out         : out   std_logic_vector(0 to 0);
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f0_out_valid : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_fifo
    port( data_wen              : in    std_logic_vector(3 downto 0) := (others => 'U');
          data_ren              : in    std_logic_vector(3 downto 0) := (others => 'U');
          ready_i_0             : out   std_logic_vector(3 downto 0);
          time_ren              : in    std_logic_vector(3 downto 0) := (others => 'U');
          time_wen              : in    std_logic_vector(3 downto 0) := (others => 'U');
          wdata                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          hwdata_c              : out   std_logic_vector(31 downto 0);
          time_ren_1z           : in    std_logic := 'U';
          data_ren_1z           : in    std_logic := 'U';
          un20_time_write       : in    std_logic := 'U';
          un13_time_write       : in    std_logic := 'U';
          HRESETn_c             : in    std_logic := 'U';
          lpp_waveform_fifo_VCC : in    std_logic := 'U';
          lpp_waveform_fifo_GND : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_snapshot_160_11
    port( sample_f0_wdata_95 : in    std_logic := 'U';
          sample_f0_wdata_94 : in    std_logic := 'U';
          sample_f0_wdata_93 : in    std_logic := 'U';
          sample_f0_wdata_92 : in    std_logic := 'U';
          sample_f0_wdata_91 : in    std_logic := 'U';
          sample_f0_wdata_90 : in    std_logic := 'U';
          sample_f0_wdata_89 : in    std_logic := 'U';
          sample_f0_wdata_88 : in    std_logic := 'U';
          sample_f0_wdata_87 : in    std_logic := 'U';
          sample_f0_wdata_86 : in    std_logic := 'U';
          sample_f0_wdata_85 : in    std_logic := 'U';
          sample_f0_wdata_84 : in    std_logic := 'U';
          sample_f0_wdata_83 : in    std_logic := 'U';
          sample_f0_wdata_82 : in    std_logic := 'U';
          sample_f0_wdata_81 : in    std_logic := 'U';
          sample_f0_wdata_80 : in    std_logic := 'U';
          sample_f0_wdata_79 : in    std_logic := 'U';
          sample_f0_wdata_78 : in    std_logic := 'U';
          sample_f0_wdata_77 : in    std_logic := 'U';
          sample_f0_wdata_76 : in    std_logic := 'U';
          sample_f0_wdata_75 : in    std_logic := 'U';
          sample_f0_wdata_74 : in    std_logic := 'U';
          sample_f0_wdata_73 : in    std_logic := 'U';
          sample_f0_wdata_72 : in    std_logic := 'U';
          sample_f0_wdata_71 : in    std_logic := 'U';
          sample_f0_wdata_70 : in    std_logic := 'U';
          sample_f0_wdata_69 : in    std_logic := 'U';
          sample_f0_wdata_68 : in    std_logic := 'U';
          sample_f0_wdata_67 : in    std_logic := 'U';
          sample_f0_wdata_66 : in    std_logic := 'U';
          sample_f0_wdata_65 : in    std_logic := 'U';
          sample_f0_wdata_64 : in    std_logic := 'U';
          sample_f0_wdata_63 : in    std_logic := 'U';
          sample_f0_wdata_62 : in    std_logic := 'U';
          sample_f0_wdata_61 : in    std_logic := 'U';
          sample_f0_wdata_60 : in    std_logic := 'U';
          sample_f0_wdata_59 : in    std_logic := 'U';
          sample_f0_wdata_58 : in    std_logic := 'U';
          sample_f0_wdata_57 : in    std_logic := 'U';
          sample_f0_wdata_56 : in    std_logic := 'U';
          sample_f0_wdata_55 : in    std_logic := 'U';
          sample_f0_wdata_54 : in    std_logic := 'U';
          sample_f0_wdata_53 : in    std_logic := 'U';
          sample_f0_wdata_52 : in    std_logic := 'U';
          sample_f0_wdata_51 : in    std_logic := 'U';
          sample_f0_wdata_50 : in    std_logic := 'U';
          sample_f0_wdata_49 : in    std_logic := 'U';
          sample_f0_wdata_48 : in    std_logic := 'U';
          sample_f0_wdata_15 : in    std_logic := 'U';
          sample_f0_wdata_14 : in    std_logic := 'U';
          sample_f0_wdata_13 : in    std_logic := 'U';
          sample_f0_wdata_12 : in    std_logic := 'U';
          sample_f0_wdata_11 : in    std_logic := 'U';
          sample_f0_wdata_10 : in    std_logic := 'U';
          sample_f0_wdata_9  : in    std_logic := 'U';
          sample_f0_wdata_8  : in    std_logic := 'U';
          sample_f0_wdata_7  : in    std_logic := 'U';
          sample_f0_wdata_6  : in    std_logic := 'U';
          sample_f0_wdata_5  : in    std_logic := 'U';
          sample_f0_wdata_4  : in    std_logic := 'U';
          sample_f0_wdata_3  : in    std_logic := 'U';
          sample_f0_wdata_2  : in    std_logic := 'U';
          sample_f0_wdata_1  : in    std_logic := 'U';
          sample_f0_wdata_0  : in    std_logic := 'U';
          data_f0_out        : out   std_logic_vector(159 downto 64);
          nb_snapshot_param  : in    std_logic_vector(10 downto 0) := (others => 'U');
          sample_f0_37       : in    std_logic := 'U';
          sample_f0_5        : in    std_logic := 'U';
          sample_f0_38       : in    std_logic := 'U';
          sample_f0_6        : in    std_logic := 'U';
          sample_f0_39       : in    std_logic := 'U';
          sample_f0_7        : in    std_logic := 'U';
          sample_f0_40       : in    std_logic := 'U';
          sample_f0_8        : in    std_logic := 'U';
          sample_f0_41       : in    std_logic := 'U';
          sample_f0_9        : in    std_logic := 'U';
          sample_f0_42       : in    std_logic := 'U';
          sample_f0_10       : in    std_logic := 'U';
          sample_f0_43       : in    std_logic := 'U';
          sample_f0_11       : in    std_logic := 'U';
          sample_f0_61       : in    std_logic := 'U';
          sample_f0_62       : in    std_logic := 'U';
          sample_f0_63       : in    std_logic := 'U';
          sample_f0_32       : in    std_logic := 'U';
          sample_f0_0        : in    std_logic := 'U';
          sample_f0_33       : in    std_logic := 'U';
          sample_f0_1        : in    std_logic := 'U';
          sample_f0_34       : in    std_logic := 'U';
          sample_f0_2        : in    std_logic := 'U';
          sample_f0_35       : in    std_logic := 'U';
          sample_f0_3        : in    std_logic := 'U';
          sample_f0_36       : in    std_logic := 'U';
          sample_f0_4        : in    std_logic := 'U';
          sample_f0_48       : in    std_logic := 'U';
          sample_f0_49       : in    std_logic := 'U';
          sample_f0_50       : in    std_logic := 'U';
          sample_f0_51       : in    std_logic := 'U';
          sample_f0_52       : in    std_logic := 'U';
          sample_f0_53       : in    std_logic := 'U';
          sample_f0_54       : in    std_logic := 'U';
          sample_f0_55       : in    std_logic := 'U';
          sample_f0_56       : in    std_logic := 'U';
          sample_f0_57       : in    std_logic := 'U';
          sample_f0_58       : in    std_logic := 'U';
          sample_f0_59       : in    std_logic := 'U';
          sample_f0_60       : in    std_logic := 'U';
          sample_f0_44       : in    std_logic := 'U';
          sample_f0_12       : in    std_logic := 'U';
          sample_f0_45       : in    std_logic := 'U';
          sample_f0_13       : in    std_logic := 'U';
          sample_f0_46       : in    std_logic := 'U';
          sample_f0_14       : in    std_logic := 'U';
          sample_f0_47       : in    std_logic := 'U';
          sample_f0_15       : in    std_logic := 'U';
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          data_f0_out_valid  : out   std_logic;
          enable_f0          : in    std_logic := 'U';
          data_shaping_R0    : in    std_logic := 'U';
          data_shaping_R0_0  : in    std_logic := 'U';
          start_snapshot_f0  : in    std_logic := 'U';
          sample_f0_val_0    : in    std_logic := 'U';
          burst_f0           : in    std_logic := 'U'
        );
  end component;

  component 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1
    port( sample_f2_wdata   : in    std_logic_vector(95 downto 0) := (others => 'U');
          data_f2_out       : out   std_logic_vector(159 downto 64);
          nb_snapshot_param : in    std_logic_vector(0 to 0) := (others => 'U');
          HRESETn_c         : in    std_logic := 'U';
          HCLK_c            : in    std_logic := 'U';
          data_f2_out_valid : out   std_logic;
          I_13_20           : in    std_logic := 'U';
          I_9_20            : in    std_logic := 'U';
          I_5_20            : in    std_logic := 'U';
          I_38_4            : in    std_logic := 'U';
          I_31_5            : in    std_logic := 'U';
          N_4               : in    std_logic := 'U';
          I_45_4            : in    std_logic := 'U';
          I_56_4            : in    std_logic := 'U';
          I_52_4            : in    std_logic := 'U';
          I_24_4            : in    std_logic := 'U';
          I_20_12           : in    std_logic := 'U';
          enable_f2         : in    std_logic := 'U';
          burst_f2          : in    std_logic := 'U';
          start_snapshot_f2 : in    std_logic := 'U';
          sample_f2_val     : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_dma
    port( addr_data_f0       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f1       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f2       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f3       : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full        : out   std_logic_vector(3 downto 0);
          status_full_err    : out   std_logic_vector(3 downto 0);
          nb_burst_available : in    std_logic_vector(10 downto 0) := (others => 'U');
          haddr_c            : out   std_logic_vector(31 downto 0);
          AHB_Master_In_c_3  : in    std_logic := 'U';
          AHB_Master_In_c_0  : in    std_logic := 'U';
          AHB_Master_In_c_4  : in    std_logic := 'U';
          AHB_Master_In_c_5  : in    std_logic := 'U';
          hsize_c            : out   std_logic_vector(1 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          hburst_c           : out   std_logic_vector(2 downto 0);
          status_full_ack    : in    std_logic_vector(3 downto 0) := (others => 'U');
          ready_i_0          : in    std_logic_vector(3 downto 0) := (others => 'U');
          data_ren           : out   std_logic_vector(3 downto 0);
          time_ren           : out   std_logic_vector(3 downto 0);
          time_ren_1z        : out   std_logic;
          data_ren_1z        : out   std_logic;
          N_43               : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          hwrite_c           : out   std_logic;
          un20_time_write    : out   std_logic;
          un13_time_write    : out   std_logic;
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U'
        );
  end component;

  component lpp_waveform_fifo_arbiter
    port( wdata       : out   std_logic_vector(31 downto 0);
          data_wen    : out   std_logic_vector(3 downto 0);
          valid_ack   : out   std_logic_vector(3 downto 0);
          time_wen    : out   std_logic_vector(3 downto 0);
          data_f3_out : in    std_logic_vector(159 downto 64) := (others => 'U');
          data_f2_out : in    std_logic_vector(159 downto 64) := (others => 'U');
          data_f1_out : in    std_logic_vector(159 downto 64) := (others => 'U');
          data_f0_out : in    std_logic_vector(159 downto 64) := (others => 'U');
          valid_out_i : in    std_logic_vector(1 to 1) := (others => 'U');
          ready_i_0   : in    std_logic_vector(3 downto 0) := (others => 'U');
          valid_out_3 : in    std_logic := 'U';
          valid_out_2 : in    std_logic := 'U';
          valid_out_0 : in    std_logic := 'U';
          HRESETn_c   : in    std_logic := 'U';
          HCLK_c      : in    std_logic := 'U'
        );
  end component;

    signal N_45, N_37, \DWACT_FINC_E[0]\, N_14, 
        \DWACT_FINC_E[4]\, N_4, \DWACT_FINC_E[6]\, 
        \DWACT_FINC_E[2]\, \DWACT_FINC_E[5]\, I_56_4, N_11, 
        I_52_4, \DWACT_FINC_E[3]\, I_45_4, N_19, I_38_4, N_24, 
        I_31_5, N_29, \DWACT_FINC_E[1]\, I_24_4, N_34, I_20_12, 
        I_13_20, N_42, I_9_20, I_5_20, start_snapshot_f2, 
        start_snapshot_f1, start_snapshot_f0, \data_f0_out[64]\, 
        \data_f0_out[65]\, \data_f0_out[66]\, \data_f0_out[67]\, 
        \data_f0_out[68]\, \data_f0_out[69]\, \data_f0_out[70]\, 
        \data_f0_out[71]\, \data_f0_out[72]\, \data_f0_out[73]\, 
        \data_f0_out[74]\, \data_f0_out[75]\, \data_f0_out[76]\, 
        \data_f0_out[77]\, \data_f0_out[78]\, \data_f0_out[79]\, 
        \data_f0_out[80]\, \data_f0_out[81]\, \data_f0_out[82]\, 
        \data_f0_out[83]\, \data_f0_out[84]\, \data_f0_out[85]\, 
        \data_f0_out[86]\, \data_f0_out[87]\, \data_f0_out[88]\, 
        \data_f0_out[89]\, \data_f0_out[90]\, \data_f0_out[91]\, 
        \data_f0_out[92]\, \data_f0_out[93]\, \data_f0_out[94]\, 
        \data_f0_out[95]\, \data_f0_out[96]\, \data_f0_out[97]\, 
        \data_f0_out[98]\, \data_f0_out[99]\, \data_f0_out[100]\, 
        \data_f0_out[101]\, \data_f0_out[102]\, 
        \data_f0_out[103]\, \data_f0_out[104]\, 
        \data_f0_out[105]\, \data_f0_out[106]\, 
        \data_f0_out[107]\, \data_f0_out[108]\, 
        \data_f0_out[109]\, \data_f0_out[110]\, 
        \data_f0_out[111]\, \data_f0_out[112]\, 
        \data_f0_out[113]\, \data_f0_out[114]\, 
        \data_f0_out[115]\, \data_f0_out[116]\, 
        \data_f0_out[117]\, \data_f0_out[118]\, 
        \data_f0_out[119]\, \data_f0_out[120]\, 
        \data_f0_out[121]\, \data_f0_out[122]\, 
        \data_f0_out[123]\, \data_f0_out[124]\, 
        \data_f0_out[125]\, \data_f0_out[126]\, 
        \data_f0_out[127]\, \data_f0_out[128]\, 
        \data_f0_out[129]\, \data_f0_out[130]\, 
        \data_f0_out[131]\, \data_f0_out[132]\, 
        \data_f0_out[133]\, \data_f0_out[134]\, 
        \data_f0_out[135]\, \data_f0_out[136]\, 
        \data_f0_out[137]\, \data_f0_out[138]\, 
        \data_f0_out[139]\, \data_f0_out[140]\, 
        \data_f0_out[141]\, \data_f0_out[142]\, 
        \data_f0_out[143]\, \data_f0_out[144]\, 
        \data_f0_out[145]\, \data_f0_out[146]\, 
        \data_f0_out[147]\, \data_f0_out[148]\, 
        \data_f0_out[149]\, \data_f0_out[150]\, 
        \data_f0_out[151]\, \data_f0_out[152]\, 
        \data_f0_out[153]\, \data_f0_out[154]\, 
        \data_f0_out[155]\, \data_f0_out[156]\, 
        \data_f0_out[157]\, \data_f0_out[158]\, 
        \data_f0_out[159]\, data_f0_out_valid, \data_f1_out[64]\, 
        \data_f1_out[65]\, \data_f1_out[66]\, \data_f1_out[67]\, 
        \data_f1_out[68]\, \data_f1_out[69]\, \data_f1_out[70]\, 
        \data_f1_out[71]\, \data_f1_out[72]\, \data_f1_out[73]\, 
        \data_f1_out[74]\, \data_f1_out[75]\, \data_f1_out[76]\, 
        \data_f1_out[77]\, \data_f1_out[78]\, \data_f1_out[79]\, 
        \data_f1_out[80]\, \data_f1_out[81]\, \data_f1_out[82]\, 
        \data_f1_out[83]\, \data_f1_out[84]\, \data_f1_out[85]\, 
        \data_f1_out[86]\, \data_f1_out[87]\, \data_f1_out[88]\, 
        \data_f1_out[89]\, \data_f1_out[90]\, \data_f1_out[91]\, 
        \data_f1_out[92]\, \data_f1_out[93]\, \data_f1_out[94]\, 
        \data_f1_out[95]\, \data_f1_out[96]\, \data_f1_out[97]\, 
        \data_f1_out[98]\, \data_f1_out[99]\, \data_f1_out[100]\, 
        \data_f1_out[101]\, \data_f1_out[102]\, 
        \data_f1_out[103]\, \data_f1_out[104]\, 
        \data_f1_out[105]\, \data_f1_out[106]\, 
        \data_f1_out[107]\, \data_f1_out[108]\, 
        \data_f1_out[109]\, \data_f1_out[110]\, 
        \data_f1_out[111]\, \data_f1_out[112]\, 
        \data_f1_out[113]\, \data_f1_out[114]\, 
        \data_f1_out[115]\, \data_f1_out[116]\, 
        \data_f1_out[117]\, \data_f1_out[118]\, 
        \data_f1_out[119]\, \data_f1_out[120]\, 
        \data_f1_out[121]\, \data_f1_out[122]\, 
        \data_f1_out[123]\, \data_f1_out[124]\, 
        \data_f1_out[125]\, \data_f1_out[126]\, 
        \data_f1_out[127]\, \data_f1_out[128]\, 
        \data_f1_out[129]\, \data_f1_out[130]\, 
        \data_f1_out[131]\, \data_f1_out[132]\, 
        \data_f1_out[133]\, \data_f1_out[134]\, 
        \data_f1_out[135]\, \data_f1_out[136]\, 
        \data_f1_out[137]\, \data_f1_out[138]\, 
        \data_f1_out[139]\, \data_f1_out[140]\, 
        \data_f1_out[141]\, \data_f1_out[142]\, 
        \data_f1_out[143]\, \data_f1_out[144]\, 
        \data_f1_out[145]\, \data_f1_out[146]\, 
        \data_f1_out[147]\, \data_f1_out[148]\, 
        \data_f1_out[149]\, \data_f1_out[150]\, 
        \data_f1_out[151]\, \data_f1_out[152]\, 
        \data_f1_out[153]\, \data_f1_out[154]\, 
        \data_f1_out[155]\, \data_f1_out[156]\, 
        \data_f1_out[157]\, \data_f1_out[158]\, 
        \data_f1_out[159]\, data_f1_out_valid, \data_f2_out[64]\, 
        \data_f2_out[65]\, \data_f2_out[66]\, \data_f2_out[67]\, 
        \data_f2_out[68]\, \data_f2_out[69]\, \data_f2_out[70]\, 
        \data_f2_out[71]\, \data_f2_out[72]\, \data_f2_out[73]\, 
        \data_f2_out[74]\, \data_f2_out[75]\, \data_f2_out[76]\, 
        \data_f2_out[77]\, \data_f2_out[78]\, \data_f2_out[79]\, 
        \data_f2_out[80]\, \data_f2_out[81]\, \data_f2_out[82]\, 
        \data_f2_out[83]\, \data_f2_out[84]\, \data_f2_out[85]\, 
        \data_f2_out[86]\, \data_f2_out[87]\, \data_f2_out[88]\, 
        \data_f2_out[89]\, \data_f2_out[90]\, \data_f2_out[91]\, 
        \data_f2_out[92]\, \data_f2_out[93]\, \data_f2_out[94]\, 
        \data_f2_out[95]\, \data_f2_out[96]\, \data_f2_out[97]\, 
        \data_f2_out[98]\, \data_f2_out[99]\, \data_f2_out[100]\, 
        \data_f2_out[101]\, \data_f2_out[102]\, 
        \data_f2_out[103]\, \data_f2_out[104]\, 
        \data_f2_out[105]\, \data_f2_out[106]\, 
        \data_f2_out[107]\, \data_f2_out[108]\, 
        \data_f2_out[109]\, \data_f2_out[110]\, 
        \data_f2_out[111]\, \data_f2_out[112]\, 
        \data_f2_out[113]\, \data_f2_out[114]\, 
        \data_f2_out[115]\, \data_f2_out[116]\, 
        \data_f2_out[117]\, \data_f2_out[118]\, 
        \data_f2_out[119]\, \data_f2_out[120]\, 
        \data_f2_out[121]\, \data_f2_out[122]\, 
        \data_f2_out[123]\, \data_f2_out[124]\, 
        \data_f2_out[125]\, \data_f2_out[126]\, 
        \data_f2_out[127]\, \data_f2_out[128]\, 
        \data_f2_out[129]\, \data_f2_out[130]\, 
        \data_f2_out[131]\, \data_f2_out[132]\, 
        \data_f2_out[133]\, \data_f2_out[134]\, 
        \data_f2_out[135]\, \data_f2_out[136]\, 
        \data_f2_out[137]\, \data_f2_out[138]\, 
        \data_f2_out[139]\, \data_f2_out[140]\, 
        \data_f2_out[141]\, \data_f2_out[142]\, 
        \data_f2_out[143]\, \data_f2_out[144]\, 
        \data_f2_out[145]\, \data_f2_out[146]\, 
        \data_f2_out[147]\, \data_f2_out[148]\, 
        \data_f2_out[149]\, \data_f2_out[150]\, 
        \data_f2_out[151]\, \data_f2_out[152]\, 
        \data_f2_out[153]\, \data_f2_out[154]\, 
        \data_f2_out[155]\, \data_f2_out[156]\, 
        \data_f2_out[157]\, \data_f2_out[158]\, 
        \data_f2_out[159]\, data_f2_out_valid, \data_f3_out[64]\, 
        \data_f3_out[65]\, \data_f3_out[66]\, \data_f3_out[67]\, 
        \data_f3_out[68]\, \data_f3_out[69]\, \data_f3_out[70]\, 
        \data_f3_out[71]\, \data_f3_out[72]\, \data_f3_out[73]\, 
        \data_f3_out[74]\, \data_f3_out[75]\, \data_f3_out[76]\, 
        \data_f3_out[77]\, \data_f3_out[78]\, \data_f3_out[79]\, 
        \data_f3_out[80]\, \data_f3_out[81]\, \data_f3_out[82]\, 
        \data_f3_out[83]\, \data_f3_out[84]\, \data_f3_out[85]\, 
        \data_f3_out[86]\, \data_f3_out[87]\, \data_f3_out[88]\, 
        \data_f3_out[89]\, \data_f3_out[90]\, \data_f3_out[91]\, 
        \data_f3_out[92]\, \data_f3_out[93]\, \data_f3_out[94]\, 
        \data_f3_out[95]\, \data_f3_out[96]\, \data_f3_out[97]\, 
        \data_f3_out[98]\, \data_f3_out[99]\, \data_f3_out[100]\, 
        \data_f3_out[101]\, \data_f3_out[102]\, 
        \data_f3_out[103]\, \data_f3_out[104]\, 
        \data_f3_out[105]\, \data_f3_out[106]\, 
        \data_f3_out[107]\, \data_f3_out[108]\, 
        \data_f3_out[109]\, \data_f3_out[110]\, 
        \data_f3_out[111]\, \data_f3_out[112]\, 
        \data_f3_out[113]\, \data_f3_out[114]\, 
        \data_f3_out[115]\, \data_f3_out[116]\, 
        \data_f3_out[117]\, \data_f3_out[118]\, 
        \data_f3_out[119]\, \data_f3_out[120]\, 
        \data_f3_out[121]\, \data_f3_out[122]\, 
        \data_f3_out[123]\, \data_f3_out[124]\, 
        \data_f3_out[125]\, \data_f3_out[126]\, 
        \data_f3_out[127]\, \data_f3_out[128]\, 
        \data_f3_out[129]\, \data_f3_out[130]\, 
        \data_f3_out[131]\, \data_f3_out[132]\, 
        \data_f3_out[133]\, \data_f3_out[134]\, 
        \data_f3_out[135]\, \data_f3_out[136]\, 
        \data_f3_out[137]\, \data_f3_out[138]\, 
        \data_f3_out[139]\, \data_f3_out[140]\, 
        \data_f3_out[141]\, \data_f3_out[142]\, 
        \data_f3_out[143]\, \data_f3_out[144]\, 
        \data_f3_out[145]\, \data_f3_out[146]\, 
        \data_f3_out[147]\, \data_f3_out[148]\, 
        \data_f3_out[149]\, \data_f3_out[150]\, 
        \data_f3_out[151]\, \data_f3_out[152]\, 
        \data_f3_out[153]\, \data_f3_out[154]\, 
        \data_f3_out[155]\, \data_f3_out[156]\, 
        \data_f3_out[157]\, \data_f3_out[158]\, 
        \data_f3_out[159]\, data_f3_out_valid, \valid_ack[3]\, 
        \valid_out[3]\, \valid_ack[0]\, \valid_out[0]\, 
        \valid_out_i[1]\, \valid_ack[1]\, \valid_ack[2]\, 
        \valid_out[2]\, \wdata[0]\, \wdata[1]\, \wdata[2]\, 
        \wdata[3]\, \wdata[4]\, \wdata[5]\, \wdata[6]\, 
        \wdata[7]\, \wdata[8]\, \wdata[9]\, \wdata[10]\, 
        \wdata[11]\, \wdata[12]\, \wdata[13]\, \wdata[14]\, 
        \wdata[15]\, \wdata[16]\, \wdata[17]\, \wdata[18]\, 
        \wdata[19]\, \wdata[20]\, \wdata[21]\, \wdata[22]\, 
        \wdata[23]\, \wdata[24]\, \wdata[25]\, \wdata[26]\, 
        \wdata[27]\, \wdata[28]\, \wdata[29]\, \wdata[30]\, 
        \wdata[31]\, \data_wen[0]\, \data_wen[1]\, \data_wen[2]\, 
        \data_wen[3]\, \time_wen[0]\, \time_wen[1]\, 
        \time_wen[2]\, \time_wen[3]\, \ready_i_0[0]\, 
        \ready_i_0[1]\, \ready_i_0[2]\, \ready_i_0[3]\, 
        \data_ren[0]\, \data_ren[1]\, \data_ren[2]\, 
        \data_ren[3]\, \time_ren[0]\, \time_ren[1]\, 
        \time_ren[2]\, \time_ren[3]\, time_ren, data_ren, 
        un20_time_write, un13_time_write, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

    for all : lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1
	Use entity work.
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1(DEF_ARCH);
    for all : lpp_waveform_snapshot_controler
	Use entity work.lpp_waveform_snapshot_controler(DEF_ARCH);
    for all : \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\
	Use entity work.
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\(DEF_ARCH);
    for all : \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\
	Use entity work.
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\(DEF_ARCH);
    for all : lpp_waveform_burst
	Use entity work.lpp_waveform_burst(DEF_ARCH);
    for all : \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\
	Use entity work.
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\(DEF_ARCH);
    for all : \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\
	Use entity work.
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\(DEF_ARCH);
    for all : lpp_waveform_fifo
	Use entity work.lpp_waveform_fifo(DEF_ARCH);
    for all : lpp_waveform_snapshot_160_11
	Use entity work.lpp_waveform_snapshot_160_11(DEF_ARCH);
    for all : lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1
	Use entity work.
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1(DEF_ARCH);
    for all : lpp_waveform_dma
	Use entity work.lpp_waveform_dma(DEF_ARCH);
    for all : lpp_waveform_fifo_arbiter
	Use entity work.lpp_waveform_fifo_arbiter(DEF_ARCH);
begin 


    un7_nb_snapshot_param_more_one_I_45 : XOR2
      port map(A => N_19, B => nb_snapshot_param(8), Y => I_45_4);
    
    un7_nb_snapshot_param_more_one_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => nb_snapshot_param(6), Y => N_24);
    
    un7_nb_snapshot_param_more_one_I_16 : AND3
      port map(A => nb_snapshot_param(0), B => 
        nb_snapshot_param(1), C => nb_snapshot_param(2), Y => 
        \DWACT_FINC_E[0]\);
    
    lpp_waveform_snapshot_f1 : 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1
      port map(sample_f1_wdata_95 => sample_f1_wdata_95, 
        sample_f1_wdata_94 => sample_f1_wdata_94, 
        sample_f1_wdata_93 => sample_f1_wdata_93, 
        sample_f1_wdata_92 => sample_f1_wdata_92, 
        sample_f1_wdata_91 => sample_f1_wdata_91, 
        sample_f1_wdata_90 => sample_f1_wdata_90, 
        sample_f1_wdata_89 => sample_f1_wdata_89, 
        sample_f1_wdata_88 => sample_f1_wdata_88, 
        sample_f1_wdata_87 => sample_f1_wdata_87, 
        sample_f1_wdata_86 => sample_f1_wdata_86, 
        sample_f1_wdata_85 => sample_f1_wdata_85, 
        sample_f1_wdata_84 => sample_f1_wdata_84, 
        sample_f1_wdata_83 => sample_f1_wdata_83, 
        sample_f1_wdata_82 => sample_f1_wdata_82, 
        sample_f1_wdata_81 => sample_f1_wdata_81, 
        sample_f1_wdata_80 => sample_f1_wdata_80, 
        sample_f1_wdata_79 => sample_f1_wdata_79, 
        sample_f1_wdata_78 => sample_f1_wdata_78, 
        sample_f1_wdata_77 => sample_f1_wdata_77, 
        sample_f1_wdata_76 => sample_f1_wdata_76, 
        sample_f1_wdata_75 => sample_f1_wdata_75, 
        sample_f1_wdata_74 => sample_f1_wdata_74, 
        sample_f1_wdata_73 => sample_f1_wdata_73, 
        sample_f1_wdata_72 => sample_f1_wdata_72, 
        sample_f1_wdata_71 => sample_f1_wdata_71, 
        sample_f1_wdata_70 => sample_f1_wdata_70, 
        sample_f1_wdata_69 => sample_f1_wdata_69, 
        sample_f1_wdata_68 => sample_f1_wdata_68, 
        sample_f1_wdata_67 => sample_f1_wdata_67, 
        sample_f1_wdata_66 => sample_f1_wdata_66, 
        sample_f1_wdata_65 => sample_f1_wdata_65, 
        sample_f1_wdata_64 => sample_f1_wdata_64, 
        sample_f1_wdata_63 => sample_f1_wdata_63, 
        sample_f1_wdata_62 => sample_f1_wdata_62, 
        sample_f1_wdata_61 => sample_f1_wdata_61, 
        sample_f1_wdata_60 => sample_f1_wdata_60, 
        sample_f1_wdata_59 => sample_f1_wdata_59, 
        sample_f1_wdata_58 => sample_f1_wdata_58, 
        sample_f1_wdata_57 => sample_f1_wdata_57, 
        sample_f1_wdata_56 => sample_f1_wdata_56, 
        sample_f1_wdata_55 => sample_f1_wdata_55, 
        sample_f1_wdata_54 => sample_f1_wdata_54, 
        sample_f1_wdata_53 => sample_f1_wdata_53, 
        sample_f1_wdata_52 => sample_f1_wdata_52, 
        sample_f1_wdata_51 => sample_f1_wdata_51, 
        sample_f1_wdata_50 => sample_f1_wdata_50, 
        sample_f1_wdata_49 => sample_f1_wdata_49, 
        sample_f1_wdata_48 => sample_f1_wdata_48, 
        sample_f1_wdata_15 => sample_f1_wdata_15, 
        sample_f1_wdata_14 => sample_f1_wdata_14, 
        sample_f1_wdata_13 => sample_f1_wdata_13, 
        sample_f1_wdata_12 => sample_f1_wdata_12, 
        sample_f1_wdata_11 => sample_f1_wdata_11, 
        sample_f1_wdata_10 => sample_f1_wdata_10, 
        sample_f1_wdata_9 => sample_f1_wdata_9, sample_f1_wdata_8
         => sample_f1_wdata_8, sample_f1_wdata_7 => 
        sample_f1_wdata_7, sample_f1_wdata_6 => sample_f1_wdata_6, 
        sample_f1_wdata_5 => sample_f1_wdata_5, sample_f1_wdata_4
         => sample_f1_wdata_4, sample_f1_wdata_3 => 
        sample_f1_wdata_3, sample_f1_wdata_2 => sample_f1_wdata_2, 
        sample_f1_wdata_1 => sample_f1_wdata_1, sample_f1_wdata_0
         => sample_f1_wdata_0, data_f1_out(159) => 
        \data_f1_out[159]\, data_f1_out(158) => 
        \data_f1_out[158]\, data_f1_out(157) => 
        \data_f1_out[157]\, data_f1_out(156) => 
        \data_f1_out[156]\, data_f1_out(155) => 
        \data_f1_out[155]\, data_f1_out(154) => 
        \data_f1_out[154]\, data_f1_out(153) => 
        \data_f1_out[153]\, data_f1_out(152) => 
        \data_f1_out[152]\, data_f1_out(151) => 
        \data_f1_out[151]\, data_f1_out(150) => 
        \data_f1_out[150]\, data_f1_out(149) => 
        \data_f1_out[149]\, data_f1_out(148) => 
        \data_f1_out[148]\, data_f1_out(147) => 
        \data_f1_out[147]\, data_f1_out(146) => 
        \data_f1_out[146]\, data_f1_out(145) => 
        \data_f1_out[145]\, data_f1_out(144) => 
        \data_f1_out[144]\, data_f1_out(143) => 
        \data_f1_out[143]\, data_f1_out(142) => 
        \data_f1_out[142]\, data_f1_out(141) => 
        \data_f1_out[141]\, data_f1_out(140) => 
        \data_f1_out[140]\, data_f1_out(139) => 
        \data_f1_out[139]\, data_f1_out(138) => 
        \data_f1_out[138]\, data_f1_out(137) => 
        \data_f1_out[137]\, data_f1_out(136) => 
        \data_f1_out[136]\, data_f1_out(135) => 
        \data_f1_out[135]\, data_f1_out(134) => 
        \data_f1_out[134]\, data_f1_out(133) => 
        \data_f1_out[133]\, data_f1_out(132) => 
        \data_f1_out[132]\, data_f1_out(131) => 
        \data_f1_out[131]\, data_f1_out(130) => 
        \data_f1_out[130]\, data_f1_out(129) => 
        \data_f1_out[129]\, data_f1_out(128) => 
        \data_f1_out[128]\, data_f1_out(127) => 
        \data_f1_out[127]\, data_f1_out(126) => 
        \data_f1_out[126]\, data_f1_out(125) => 
        \data_f1_out[125]\, data_f1_out(124) => 
        \data_f1_out[124]\, data_f1_out(123) => 
        \data_f1_out[123]\, data_f1_out(122) => 
        \data_f1_out[122]\, data_f1_out(121) => 
        \data_f1_out[121]\, data_f1_out(120) => 
        \data_f1_out[120]\, data_f1_out(119) => 
        \data_f1_out[119]\, data_f1_out(118) => 
        \data_f1_out[118]\, data_f1_out(117) => 
        \data_f1_out[117]\, data_f1_out(116) => 
        \data_f1_out[116]\, data_f1_out(115) => 
        \data_f1_out[115]\, data_f1_out(114) => 
        \data_f1_out[114]\, data_f1_out(113) => 
        \data_f1_out[113]\, data_f1_out(112) => 
        \data_f1_out[112]\, data_f1_out(111) => 
        \data_f1_out[111]\, data_f1_out(110) => 
        \data_f1_out[110]\, data_f1_out(109) => 
        \data_f1_out[109]\, data_f1_out(108) => 
        \data_f1_out[108]\, data_f1_out(107) => 
        \data_f1_out[107]\, data_f1_out(106) => 
        \data_f1_out[106]\, data_f1_out(105) => 
        \data_f1_out[105]\, data_f1_out(104) => 
        \data_f1_out[104]\, data_f1_out(103) => 
        \data_f1_out[103]\, data_f1_out(102) => 
        \data_f1_out[102]\, data_f1_out(101) => 
        \data_f1_out[101]\, data_f1_out(100) => 
        \data_f1_out[100]\, data_f1_out(99) => \data_f1_out[99]\, 
        data_f1_out(98) => \data_f1_out[98]\, data_f1_out(97) => 
        \data_f1_out[97]\, data_f1_out(96) => \data_f1_out[96]\, 
        data_f1_out(95) => \data_f1_out[95]\, data_f1_out(94) => 
        \data_f1_out[94]\, data_f1_out(93) => \data_f1_out[93]\, 
        data_f1_out(92) => \data_f1_out[92]\, data_f1_out(91) => 
        \data_f1_out[91]\, data_f1_out(90) => \data_f1_out[90]\, 
        data_f1_out(89) => \data_f1_out[89]\, data_f1_out(88) => 
        \data_f1_out[88]\, data_f1_out(87) => \data_f1_out[87]\, 
        data_f1_out(86) => \data_f1_out[86]\, data_f1_out(85) => 
        \data_f1_out[85]\, data_f1_out(84) => \data_f1_out[84]\, 
        data_f1_out(83) => \data_f1_out[83]\, data_f1_out(82) => 
        \data_f1_out[82]\, data_f1_out(81) => \data_f1_out[81]\, 
        data_f1_out(80) => \data_f1_out[80]\, data_f1_out(79) => 
        \data_f1_out[79]\, data_f1_out(78) => \data_f1_out[78]\, 
        data_f1_out(77) => \data_f1_out[77]\, data_f1_out(76) => 
        \data_f1_out[76]\, data_f1_out(75) => \data_f1_out[75]\, 
        data_f1_out(74) => \data_f1_out[74]\, data_f1_out(73) => 
        \data_f1_out[73]\, data_f1_out(72) => \data_f1_out[72]\, 
        data_f1_out(71) => \data_f1_out[71]\, data_f1_out(70) => 
        \data_f1_out[70]\, data_f1_out(69) => \data_f1_out[69]\, 
        data_f1_out(68) => \data_f1_out[68]\, data_f1_out(67) => 
        \data_f1_out[67]\, data_f1_out(66) => \data_f1_out[66]\, 
        data_f1_out(65) => \data_f1_out[65]\, data_f1_out(64) => 
        \data_f1_out[64]\, nb_snapshot_param(0) => 
        nb_snapshot_param(0), sample_f1_37 => sample_f1_37, 
        sample_f1_5 => sample_f1_5, sample_f1_38 => sample_f1_38, 
        sample_f1_6 => sample_f1_6, sample_f1_39 => sample_f1_39, 
        sample_f1_7 => sample_f1_7, sample_f1_40 => sample_f1_40, 
        sample_f1_8 => sample_f1_8, sample_f1_41 => sample_f1_41, 
        sample_f1_9 => sample_f1_9, sample_f1_42 => sample_f1_42, 
        sample_f1_10 => sample_f1_10, sample_f1_43 => 
        sample_f1_43, sample_f1_11 => sample_f1_11, sample_f1_61
         => sample_f1_61, sample_f1_62 => sample_f1_62, 
        sample_f1_63 => sample_f1_63, sample_f1_32 => 
        sample_f1_32, sample_f1_0 => sample_f1_0, sample_f1_33
         => sample_f1_33, sample_f1_1 => sample_f1_1, 
        sample_f1_34 => sample_f1_34, sample_f1_2 => sample_f1_2, 
        sample_f1_35 => sample_f1_35, sample_f1_3 => sample_f1_3, 
        sample_f1_36 => sample_f1_36, sample_f1_4 => sample_f1_4, 
        sample_f1_48 => sample_f1_48, sample_f1_49 => 
        sample_f1_49, sample_f1_50 => sample_f1_50, sample_f1_51
         => sample_f1_51, sample_f1_52 => sample_f1_52, 
        sample_f1_53 => sample_f1_53, sample_f1_54 => 
        sample_f1_54, sample_f1_55 => sample_f1_55, sample_f1_56
         => sample_f1_56, sample_f1_57 => sample_f1_57, 
        sample_f1_58 => sample_f1_58, sample_f1_59 => 
        sample_f1_59, sample_f1_60 => sample_f1_60, sample_f1_44
         => sample_f1_44, sample_f1_12 => sample_f1_12, 
        sample_f1_45 => sample_f1_45, sample_f1_13 => 
        sample_f1_13, sample_f1_46 => sample_f1_46, sample_f1_14
         => sample_f1_14, sample_f1_47 => sample_f1_47, 
        sample_f1_15 => sample_f1_15, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, data_f1_out_valid => data_f1_out_valid, 
        N_4 => N_4, I_38_4 => I_38_4, I_24_4 => I_24_4, I_20_12
         => I_20_12, I_13_20 => I_13_20, I_45_4 => I_45_4, I_9_20
         => I_9_20, I_5_20 => I_5_20, I_52_4 => I_52_4, 
        data_shaping_R1 => data_shaping_R1, data_shaping_R1_0 => 
        data_shaping_R1_0, I_56_4 => I_56_4, I_31_5 => I_31_5, 
        enable_f1 => enable_f1, burst_f1 => burst_f1, 
        sample_f1_val_0 => sample_f1_val_0, start_snapshot_f1 => 
        start_snapshot_f1);
    
    lpp_waveform_snapshot_controler_1 : 
        lpp_waveform_snapshot_controler
      port map(delta_f2_f0(9) => delta_f2_f0(9), delta_f2_f0(8)
         => delta_f2_f0(8), delta_f2_f0(7) => delta_f2_f0(7), 
        delta_f2_f0(6) => delta_f2_f0(6), delta_f2_f0(5) => 
        delta_f2_f0(5), delta_f2_f0(4) => delta_f2_f0(4), 
        delta_f2_f0(3) => delta_f2_f0(3), delta_f2_f0(2) => 
        delta_f2_f0(2), delta_f2_f0(1) => delta_f2_f0(1), 
        delta_f2_f0(0) => delta_f2_f0(0), delta_snapshot(15) => 
        delta_snapshot(15), delta_snapshot(14) => 
        delta_snapshot(14), delta_snapshot(13) => 
        delta_snapshot(13), delta_snapshot(12) => 
        delta_snapshot(12), delta_snapshot(11) => 
        delta_snapshot(11), delta_snapshot(10) => 
        delta_snapshot(10), delta_snapshot(9) => 
        delta_snapshot(9), delta_snapshot(8) => delta_snapshot(8), 
        delta_snapshot(7) => delta_snapshot(7), delta_snapshot(6)
         => delta_snapshot(6), delta_snapshot(5) => 
        delta_snapshot(5), delta_snapshot(4) => delta_snapshot(4), 
        delta_snapshot(3) => delta_snapshot(3), delta_snapshot(2)
         => delta_snapshot(2), delta_snapshot(1) => 
        delta_snapshot(1), delta_snapshot(0) => delta_snapshot(0), 
        delta_f2_f1(9) => delta_f2_f1(9), delta_f2_f1(8) => 
        delta_f2_f1(8), delta_f2_f1(7) => delta_f2_f1(7), 
        delta_f2_f1(6) => delta_f2_f1(6), delta_f2_f1(5) => 
        delta_f2_f1(5), delta_f2_f1(4) => delta_f2_f1(4), 
        delta_f2_f1(3) => delta_f2_f1(3), delta_f2_f1(2) => 
        delta_f2_f1(2), delta_f2_f1(1) => delta_f2_f1(1), 
        delta_f2_f1(0) => delta_f2_f1(0), start_snapshot_f2 => 
        start_snapshot_f2, start_snapshot_f1 => start_snapshot_f1, 
        start_snapshot_f0 => start_snapshot_f0, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, sample_f0_val_0 => 
        sample_f0_val_0, sample_f2_val => sample_f2_val, 
        coarse_time_0_c => coarse_time_0_c);
    
    un7_nb_snapshot_param_more_one_I_20 : XOR2
      port map(A => N_37, B => nb_snapshot_param(4), Y => I_20_12);
    
    \all_input_valid.3.lpp_waveform_dma_gen_valid_I\ : 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I\
      port map(status_new_err(3) => status_new_err(3), 
        valid_ack(3) => \valid_ack[3]\, valid_out(3) => 
        \valid_out[3]\, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, 
        data_f3_out_valid => data_f3_out_valid);
    
    un7_nb_snapshot_param_more_one_I_52 : XOR2
      port map(A => N_14, B => nb_snapshot_param(9), Y => I_52_4);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un7_nb_snapshot_param_more_one_I_62 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[6]\);
    
    un7_nb_snapshot_param_more_one_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => nb_snapshot_param(3), 
        C => nb_snapshot_param(4), Y => N_34);
    
    un7_nb_snapshot_param_more_one_I_56 : XOR2
      port map(A => N_11, B => nb_snapshot_param(10), Y => I_56_4);
    
    un7_nb_snapshot_param_more_one_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    un7_nb_snapshot_param_more_one_I_19 : NOR2B
      port map(A => nb_snapshot_param(3), B => \DWACT_FINC_E[0]\, 
        Y => N_37);
    
    un7_nb_snapshot_param_more_one_I_24 : XOR2
      port map(A => N_34, B => nb_snapshot_param(5), Y => I_24_4);
    
    un7_nb_snapshot_param_more_one_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_19);
    
    \all_input_valid.1.lpp_waveform_dma_gen_valid_I\ : 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_2\
      port map(status_new_err(1) => status_new_err(1), 
        valid_out_i(1) => \valid_out_i[1]\, valid_ack(1) => 
        \valid_ack[1]\, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, 
        data_f1_out_valid => data_f1_out_valid);
    
    un7_nb_snapshot_param_more_one_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => nb_snapshot_param(8), 
        C => nb_snapshot_param(9), Y => N_11);
    
    un7_nb_snapshot_param_more_one_I_13 : XOR2
      port map(A => N_42, B => nb_snapshot_param(3), Y => I_13_20);
    
    un7_nb_snapshot_param_more_one_I_9 : XOR2
      port map(A => N_45, B => nb_snapshot_param(2), Y => I_9_20);
    
    un7_nb_snapshot_param_more_one_I_65 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => nb_snapshot_param(9), 
        C => nb_snapshot_param(10), Y => N_4);
    
    un7_nb_snapshot_param_more_one_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => nb_snapshot_param(5), Y => N_29);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un7_nb_snapshot_param_more_one_I_59 : AND3
      port map(A => nb_snapshot_param(6), B => 
        nb_snapshot_param(7), C => nb_snapshot_param(8), Y => 
        \DWACT_FINC_E[5]\);
    
    lpp_waveform_burst_f3 : lpp_waveform_burst
      port map(sample_f3_wdata(95) => sample_f3_wdata(95), 
        sample_f3_wdata(94) => sample_f3_wdata(94), 
        sample_f3_wdata(93) => sample_f3_wdata(93), 
        sample_f3_wdata(92) => sample_f3_wdata(92), 
        sample_f3_wdata(91) => sample_f3_wdata(91), 
        sample_f3_wdata(90) => sample_f3_wdata(90), 
        sample_f3_wdata(89) => sample_f3_wdata(89), 
        sample_f3_wdata(88) => sample_f3_wdata(88), 
        sample_f3_wdata(87) => sample_f3_wdata(87), 
        sample_f3_wdata(86) => sample_f3_wdata(86), 
        sample_f3_wdata(85) => sample_f3_wdata(85), 
        sample_f3_wdata(84) => sample_f3_wdata(84), 
        sample_f3_wdata(83) => sample_f3_wdata(83), 
        sample_f3_wdata(82) => sample_f3_wdata(82), 
        sample_f3_wdata(81) => sample_f3_wdata(81), 
        sample_f3_wdata(80) => sample_f3_wdata(80), 
        sample_f3_wdata(79) => sample_f3_wdata(79), 
        sample_f3_wdata(78) => sample_f3_wdata(78), 
        sample_f3_wdata(77) => sample_f3_wdata(77), 
        sample_f3_wdata(76) => sample_f3_wdata(76), 
        sample_f3_wdata(75) => sample_f3_wdata(75), 
        sample_f3_wdata(74) => sample_f3_wdata(74), 
        sample_f3_wdata(73) => sample_f3_wdata(73), 
        sample_f3_wdata(72) => sample_f3_wdata(72), 
        sample_f3_wdata(71) => sample_f3_wdata(71), 
        sample_f3_wdata(70) => sample_f3_wdata(70), 
        sample_f3_wdata(69) => sample_f3_wdata(69), 
        sample_f3_wdata(68) => sample_f3_wdata(68), 
        sample_f3_wdata(67) => sample_f3_wdata(67), 
        sample_f3_wdata(66) => sample_f3_wdata(66), 
        sample_f3_wdata(65) => sample_f3_wdata(65), 
        sample_f3_wdata(64) => sample_f3_wdata(64), 
        sample_f3_wdata(63) => sample_f3_wdata(63), 
        sample_f3_wdata(62) => sample_f3_wdata(62), 
        sample_f3_wdata(61) => sample_f3_wdata(61), 
        sample_f3_wdata(60) => sample_f3_wdata(60), 
        sample_f3_wdata(59) => sample_f3_wdata(59), 
        sample_f3_wdata(58) => sample_f3_wdata(58), 
        sample_f3_wdata(57) => sample_f3_wdata(57), 
        sample_f3_wdata(56) => sample_f3_wdata(56), 
        sample_f3_wdata(55) => sample_f3_wdata(55), 
        sample_f3_wdata(54) => sample_f3_wdata(54), 
        sample_f3_wdata(53) => sample_f3_wdata(53), 
        sample_f3_wdata(52) => sample_f3_wdata(52), 
        sample_f3_wdata(51) => sample_f3_wdata(51), 
        sample_f3_wdata(50) => sample_f3_wdata(50), 
        sample_f3_wdata(49) => sample_f3_wdata(49), 
        sample_f3_wdata(48) => sample_f3_wdata(48), 
        sample_f3_wdata(47) => sample_f3_wdata(47), 
        sample_f3_wdata(46) => sample_f3_wdata(46), 
        sample_f3_wdata(45) => sample_f3_wdata(45), 
        sample_f3_wdata(44) => sample_f3_wdata(44), 
        sample_f3_wdata(43) => sample_f3_wdata(43), 
        sample_f3_wdata(42) => sample_f3_wdata(42), 
        sample_f3_wdata(41) => sample_f3_wdata(41), 
        sample_f3_wdata(40) => sample_f3_wdata(40), 
        sample_f3_wdata(39) => sample_f3_wdata(39), 
        sample_f3_wdata(38) => sample_f3_wdata(38), 
        sample_f3_wdata(37) => sample_f3_wdata(37), 
        sample_f3_wdata(36) => sample_f3_wdata(36), 
        sample_f3_wdata(35) => sample_f3_wdata(35), 
        sample_f3_wdata(34) => sample_f3_wdata(34), 
        sample_f3_wdata(33) => sample_f3_wdata(33), 
        sample_f3_wdata(32) => sample_f3_wdata(32), 
        sample_f3_wdata(31) => sample_f3_wdata(31), 
        sample_f3_wdata(30) => sample_f3_wdata(30), 
        sample_f3_wdata(29) => sample_f3_wdata(29), 
        sample_f3_wdata(28) => sample_f3_wdata(28), 
        sample_f3_wdata(27) => sample_f3_wdata(27), 
        sample_f3_wdata(26) => sample_f3_wdata(26), 
        sample_f3_wdata(25) => sample_f3_wdata(25), 
        sample_f3_wdata(24) => sample_f3_wdata(24), 
        sample_f3_wdata(23) => sample_f3_wdata(23), 
        sample_f3_wdata(22) => sample_f3_wdata(22), 
        sample_f3_wdata(21) => sample_f3_wdata(21), 
        sample_f3_wdata(20) => sample_f3_wdata(20), 
        sample_f3_wdata(19) => sample_f3_wdata(19), 
        sample_f3_wdata(18) => sample_f3_wdata(18), 
        sample_f3_wdata(17) => sample_f3_wdata(17), 
        sample_f3_wdata(16) => sample_f3_wdata(16), 
        sample_f3_wdata(15) => sample_f3_wdata(15), 
        sample_f3_wdata(14) => sample_f3_wdata(14), 
        sample_f3_wdata(13) => sample_f3_wdata(13), 
        sample_f3_wdata(12) => sample_f3_wdata(12), 
        sample_f3_wdata(11) => sample_f3_wdata(11), 
        sample_f3_wdata(10) => sample_f3_wdata(10), 
        sample_f3_wdata(9) => sample_f3_wdata(9), 
        sample_f3_wdata(8) => sample_f3_wdata(8), 
        sample_f3_wdata(7) => sample_f3_wdata(7), 
        sample_f3_wdata(6) => sample_f3_wdata(6), 
        sample_f3_wdata(5) => sample_f3_wdata(5), 
        sample_f3_wdata(4) => sample_f3_wdata(4), 
        sample_f3_wdata(3) => sample_f3_wdata(3), 
        sample_f3_wdata(2) => sample_f3_wdata(2), 
        sample_f3_wdata(1) => sample_f3_wdata(1), 
        sample_f3_wdata(0) => sample_f3_wdata(0), 
        data_f3_out(159) => \data_f3_out[159]\, data_f3_out(158)
         => \data_f3_out[158]\, data_f3_out(157) => 
        \data_f3_out[157]\, data_f3_out(156) => 
        \data_f3_out[156]\, data_f3_out(155) => 
        \data_f3_out[155]\, data_f3_out(154) => 
        \data_f3_out[154]\, data_f3_out(153) => 
        \data_f3_out[153]\, data_f3_out(152) => 
        \data_f3_out[152]\, data_f3_out(151) => 
        \data_f3_out[151]\, data_f3_out(150) => 
        \data_f3_out[150]\, data_f3_out(149) => 
        \data_f3_out[149]\, data_f3_out(148) => 
        \data_f3_out[148]\, data_f3_out(147) => 
        \data_f3_out[147]\, data_f3_out(146) => 
        \data_f3_out[146]\, data_f3_out(145) => 
        \data_f3_out[145]\, data_f3_out(144) => 
        \data_f3_out[144]\, data_f3_out(143) => 
        \data_f3_out[143]\, data_f3_out(142) => 
        \data_f3_out[142]\, data_f3_out(141) => 
        \data_f3_out[141]\, data_f3_out(140) => 
        \data_f3_out[140]\, data_f3_out(139) => 
        \data_f3_out[139]\, data_f3_out(138) => 
        \data_f3_out[138]\, data_f3_out(137) => 
        \data_f3_out[137]\, data_f3_out(136) => 
        \data_f3_out[136]\, data_f3_out(135) => 
        \data_f3_out[135]\, data_f3_out(134) => 
        \data_f3_out[134]\, data_f3_out(133) => 
        \data_f3_out[133]\, data_f3_out(132) => 
        \data_f3_out[132]\, data_f3_out(131) => 
        \data_f3_out[131]\, data_f3_out(130) => 
        \data_f3_out[130]\, data_f3_out(129) => 
        \data_f3_out[129]\, data_f3_out(128) => 
        \data_f3_out[128]\, data_f3_out(127) => 
        \data_f3_out[127]\, data_f3_out(126) => 
        \data_f3_out[126]\, data_f3_out(125) => 
        \data_f3_out[125]\, data_f3_out(124) => 
        \data_f3_out[124]\, data_f3_out(123) => 
        \data_f3_out[123]\, data_f3_out(122) => 
        \data_f3_out[122]\, data_f3_out(121) => 
        \data_f3_out[121]\, data_f3_out(120) => 
        \data_f3_out[120]\, data_f3_out(119) => 
        \data_f3_out[119]\, data_f3_out(118) => 
        \data_f3_out[118]\, data_f3_out(117) => 
        \data_f3_out[117]\, data_f3_out(116) => 
        \data_f3_out[116]\, data_f3_out(115) => 
        \data_f3_out[115]\, data_f3_out(114) => 
        \data_f3_out[114]\, data_f3_out(113) => 
        \data_f3_out[113]\, data_f3_out(112) => 
        \data_f3_out[112]\, data_f3_out(111) => 
        \data_f3_out[111]\, data_f3_out(110) => 
        \data_f3_out[110]\, data_f3_out(109) => 
        \data_f3_out[109]\, data_f3_out(108) => 
        \data_f3_out[108]\, data_f3_out(107) => 
        \data_f3_out[107]\, data_f3_out(106) => 
        \data_f3_out[106]\, data_f3_out(105) => 
        \data_f3_out[105]\, data_f3_out(104) => 
        \data_f3_out[104]\, data_f3_out(103) => 
        \data_f3_out[103]\, data_f3_out(102) => 
        \data_f3_out[102]\, data_f3_out(101) => 
        \data_f3_out[101]\, data_f3_out(100) => 
        \data_f3_out[100]\, data_f3_out(99) => \data_f3_out[99]\, 
        data_f3_out(98) => \data_f3_out[98]\, data_f3_out(97) => 
        \data_f3_out[97]\, data_f3_out(96) => \data_f3_out[96]\, 
        data_f3_out(95) => \data_f3_out[95]\, data_f3_out(94) => 
        \data_f3_out[94]\, data_f3_out(93) => \data_f3_out[93]\, 
        data_f3_out(92) => \data_f3_out[92]\, data_f3_out(91) => 
        \data_f3_out[91]\, data_f3_out(90) => \data_f3_out[90]\, 
        data_f3_out(89) => \data_f3_out[89]\, data_f3_out(88) => 
        \data_f3_out[88]\, data_f3_out(87) => \data_f3_out[87]\, 
        data_f3_out(86) => \data_f3_out[86]\, data_f3_out(85) => 
        \data_f3_out[85]\, data_f3_out(84) => \data_f3_out[84]\, 
        data_f3_out(83) => \data_f3_out[83]\, data_f3_out(82) => 
        \data_f3_out[82]\, data_f3_out(81) => \data_f3_out[81]\, 
        data_f3_out(80) => \data_f3_out[80]\, data_f3_out(79) => 
        \data_f3_out[79]\, data_f3_out(78) => \data_f3_out[78]\, 
        data_f3_out(77) => \data_f3_out[77]\, data_f3_out(76) => 
        \data_f3_out[76]\, data_f3_out(75) => \data_f3_out[75]\, 
        data_f3_out(74) => \data_f3_out[74]\, data_f3_out(73) => 
        \data_f3_out[73]\, data_f3_out(72) => \data_f3_out[72]\, 
        data_f3_out(71) => \data_f3_out[71]\, data_f3_out(70) => 
        \data_f3_out[70]\, data_f3_out(69) => \data_f3_out[69]\, 
        data_f3_out(68) => \data_f3_out[68]\, data_f3_out(67) => 
        \data_f3_out[67]\, data_f3_out(66) => \data_f3_out[66]\, 
        data_f3_out(65) => \data_f3_out[65]\, data_f3_out(64) => 
        \data_f3_out[64]\, HRESETn_c => HRESETn_c, HCLK_c => 
        HCLK_c, data_f3_out_valid => data_f3_out_valid, enable_f3
         => enable_f3, sample_f3_val => sample_f3_val);
    
    \all_input_valid.2.lpp_waveform_dma_gen_valid_I\ : 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_3\
      port map(status_new_err(2) => status_new_err(2), 
        valid_ack(2) => \valid_ack[2]\, valid_out(2) => 
        \valid_out[2]\, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, 
        data_f2_out_valid => data_f2_out_valid);
    
    un7_nb_snapshot_param_more_one_I_41 : AND2
      port map(A => nb_snapshot_param(6), B => 
        nb_snapshot_param(7), Y => \DWACT_FINC_E[3]\);
    
    un7_nb_snapshot_param_more_one_I_38 : XOR2
      port map(A => N_24, B => nb_snapshot_param(7), Y => I_38_4);
    
    \all_input_valid.0.lpp_waveform_dma_gen_valid_I\ : 
        \lpp_waveform_dma_gen_valid_all_input_valid.3.lpp_waveform_dma_gen_valid_I_1\
      port map(status_new_err(0) => status_new_err(0), 
        valid_ack(0) => \valid_ack[0]\, valid_out(0) => 
        \valid_out[0]\, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, 
        data_f0_out_valid => data_f0_out_valid);
    
    un7_nb_snapshot_param_more_one_I_27 : AND2
      port map(A => nb_snapshot_param(3), B => 
        nb_snapshot_param(4), Y => \DWACT_FINC_E[1]\);
    
    un7_nb_snapshot_param_more_one_I_34 : AND3
      port map(A => nb_snapshot_param(3), B => 
        nb_snapshot_param(4), C => nb_snapshot_param(5), Y => 
        \DWACT_FINC_E[2]\);
    
    un7_nb_snapshot_param_more_one_I_8 : NOR2B
      port map(A => nb_snapshot_param(1), B => 
        nb_snapshot_param(0), Y => N_45);
    
    lpp_waveform_fifo_1 : lpp_waveform_fifo
      port map(data_wen(3) => \data_wen[3]\, data_wen(2) => 
        \data_wen[2]\, data_wen(1) => \data_wen[1]\, data_wen(0)
         => \data_wen[0]\, data_ren(3) => \data_ren[3]\, 
        data_ren(2) => \data_ren[2]\, data_ren(1) => 
        \data_ren[1]\, data_ren(0) => \data_ren[0]\, ready_i_0(3)
         => \ready_i_0[3]\, ready_i_0(2) => \ready_i_0[2]\, 
        ready_i_0(1) => \ready_i_0[1]\, ready_i_0(0) => 
        \ready_i_0[0]\, time_ren(3) => \time_ren[3]\, time_ren(2)
         => \time_ren[2]\, time_ren(1) => \time_ren[1]\, 
        time_ren(0) => \time_ren[0]\, time_wen(3) => 
        \time_wen[3]\, time_wen(2) => \time_wen[2]\, time_wen(1)
         => \time_wen[1]\, time_wen(0) => \time_wen[0]\, 
        wdata(31) => \wdata[31]\, wdata(30) => \wdata[30]\, 
        wdata(29) => \wdata[29]\, wdata(28) => \wdata[28]\, 
        wdata(27) => \wdata[27]\, wdata(26) => \wdata[26]\, 
        wdata(25) => \wdata[25]\, wdata(24) => \wdata[24]\, 
        wdata(23) => \wdata[23]\, wdata(22) => \wdata[22]\, 
        wdata(21) => \wdata[21]\, wdata(20) => \wdata[20]\, 
        wdata(19) => \wdata[19]\, wdata(18) => \wdata[18]\, 
        wdata(17) => \wdata[17]\, wdata(16) => \wdata[16]\, 
        wdata(15) => \wdata[15]\, wdata(14) => \wdata[14]\, 
        wdata(13) => \wdata[13]\, wdata(12) => \wdata[12]\, 
        wdata(11) => \wdata[11]\, wdata(10) => \wdata[10]\, 
        wdata(9) => \wdata[9]\, wdata(8) => \wdata[8]\, wdata(7)
         => \wdata[7]\, wdata(6) => \wdata[6]\, wdata(5) => 
        \wdata[5]\, wdata(4) => \wdata[4]\, wdata(3) => 
        \wdata[3]\, wdata(2) => \wdata[2]\, wdata(1) => 
        \wdata[1]\, wdata(0) => \wdata[0]\, hwdata_c(31) => 
        hwdata_c(31), hwdata_c(30) => hwdata_c(30), hwdata_c(29)
         => hwdata_c(29), hwdata_c(28) => hwdata_c(28), 
        hwdata_c(27) => hwdata_c(27), hwdata_c(26) => 
        hwdata_c(26), hwdata_c(25) => hwdata_c(25), hwdata_c(24)
         => hwdata_c(24), hwdata_c(23) => hwdata_c(23), 
        hwdata_c(22) => hwdata_c(22), hwdata_c(21) => 
        hwdata_c(21), hwdata_c(20) => hwdata_c(20), hwdata_c(19)
         => hwdata_c(19), hwdata_c(18) => hwdata_c(18), 
        hwdata_c(17) => hwdata_c(17), hwdata_c(16) => 
        hwdata_c(16), hwdata_c(15) => hwdata_c(15), hwdata_c(14)
         => hwdata_c(14), hwdata_c(13) => hwdata_c(13), 
        hwdata_c(12) => hwdata_c(12), hwdata_c(11) => 
        hwdata_c(11), hwdata_c(10) => hwdata_c(10), hwdata_c(9)
         => hwdata_c(9), hwdata_c(8) => hwdata_c(8), hwdata_c(7)
         => hwdata_c(7), hwdata_c(6) => hwdata_c(6), hwdata_c(5)
         => hwdata_c(5), hwdata_c(4) => hwdata_c(4), hwdata_c(3)
         => hwdata_c(3), hwdata_c(2) => hwdata_c(2), hwdata_c(1)
         => hwdata_c(1), hwdata_c(0) => hwdata_c(0), time_ren_1z
         => time_ren, data_ren_1z => data_ren, un20_time_write
         => un20_time_write, un13_time_write => un13_time_write, 
        HRESETn_c => HRESETn_c, lpp_waveform_fifo_VCC => 
        lpp_waveform_VCC, lpp_waveform_fifo_GND => 
        lpp_waveform_GND, HCLK_c => HCLK_c);
    
    lpp_waveform_snapshot_f0 : lpp_waveform_snapshot_160_11
      port map(sample_f0_wdata_95 => sample_f0_wdata_95, 
        sample_f0_wdata_94 => sample_f0_wdata_94, 
        sample_f0_wdata_93 => sample_f0_wdata_93, 
        sample_f0_wdata_92 => sample_f0_wdata_92, 
        sample_f0_wdata_91 => sample_f0_wdata_91, 
        sample_f0_wdata_90 => sample_f0_wdata_90, 
        sample_f0_wdata_89 => sample_f0_wdata_89, 
        sample_f0_wdata_88 => sample_f0_wdata_88, 
        sample_f0_wdata_87 => sample_f0_wdata_87, 
        sample_f0_wdata_86 => sample_f0_wdata_86, 
        sample_f0_wdata_85 => sample_f0_wdata_85, 
        sample_f0_wdata_84 => sample_f0_wdata_84, 
        sample_f0_wdata_83 => sample_f0_wdata_83, 
        sample_f0_wdata_82 => sample_f0_wdata_82, 
        sample_f0_wdata_81 => sample_f0_wdata_81, 
        sample_f0_wdata_80 => sample_f0_wdata_80, 
        sample_f0_wdata_79 => sample_f0_wdata_79, 
        sample_f0_wdata_78 => sample_f0_wdata_78, 
        sample_f0_wdata_77 => sample_f0_wdata_77, 
        sample_f0_wdata_76 => sample_f0_wdata_76, 
        sample_f0_wdata_75 => sample_f0_wdata_75, 
        sample_f0_wdata_74 => sample_f0_wdata_74, 
        sample_f0_wdata_73 => sample_f0_wdata_73, 
        sample_f0_wdata_72 => sample_f0_wdata_72, 
        sample_f0_wdata_71 => sample_f0_wdata_71, 
        sample_f0_wdata_70 => sample_f0_wdata_70, 
        sample_f0_wdata_69 => sample_f0_wdata_69, 
        sample_f0_wdata_68 => sample_f0_wdata_68, 
        sample_f0_wdata_67 => sample_f0_wdata_67, 
        sample_f0_wdata_66 => sample_f0_wdata_66, 
        sample_f0_wdata_65 => sample_f0_wdata_65, 
        sample_f0_wdata_64 => sample_f0_wdata_64, 
        sample_f0_wdata_63 => sample_f0_wdata_63, 
        sample_f0_wdata_62 => sample_f0_wdata_62, 
        sample_f0_wdata_61 => sample_f0_wdata_61, 
        sample_f0_wdata_60 => sample_f0_wdata_60, 
        sample_f0_wdata_59 => sample_f0_wdata_59, 
        sample_f0_wdata_58 => sample_f0_wdata_58, 
        sample_f0_wdata_57 => sample_f0_wdata_57, 
        sample_f0_wdata_56 => sample_f0_wdata_56, 
        sample_f0_wdata_55 => sample_f0_wdata_55, 
        sample_f0_wdata_54 => sample_f0_wdata_54, 
        sample_f0_wdata_53 => sample_f0_wdata_53, 
        sample_f0_wdata_52 => sample_f0_wdata_52, 
        sample_f0_wdata_51 => sample_f0_wdata_51, 
        sample_f0_wdata_50 => sample_f0_wdata_50, 
        sample_f0_wdata_49 => sample_f0_wdata_49, 
        sample_f0_wdata_48 => sample_f0_wdata_48, 
        sample_f0_wdata_15 => sample_f0_wdata_15, 
        sample_f0_wdata_14 => sample_f0_wdata_14, 
        sample_f0_wdata_13 => sample_f0_wdata_13, 
        sample_f0_wdata_12 => sample_f0_wdata_12, 
        sample_f0_wdata_11 => sample_f0_wdata_11, 
        sample_f0_wdata_10 => sample_f0_wdata_10, 
        sample_f0_wdata_9 => sample_f0_wdata_9, sample_f0_wdata_8
         => sample_f0_wdata_8, sample_f0_wdata_7 => 
        sample_f0_wdata_7, sample_f0_wdata_6 => sample_f0_wdata_6, 
        sample_f0_wdata_5 => sample_f0_wdata_5, sample_f0_wdata_4
         => sample_f0_wdata_4, sample_f0_wdata_3 => 
        sample_f0_wdata_3, sample_f0_wdata_2 => sample_f0_wdata_2, 
        sample_f0_wdata_1 => sample_f0_wdata_1, sample_f0_wdata_0
         => sample_f0_wdata_0, data_f0_out(159) => 
        \data_f0_out[159]\, data_f0_out(158) => 
        \data_f0_out[158]\, data_f0_out(157) => 
        \data_f0_out[157]\, data_f0_out(156) => 
        \data_f0_out[156]\, data_f0_out(155) => 
        \data_f0_out[155]\, data_f0_out(154) => 
        \data_f0_out[154]\, data_f0_out(153) => 
        \data_f0_out[153]\, data_f0_out(152) => 
        \data_f0_out[152]\, data_f0_out(151) => 
        \data_f0_out[151]\, data_f0_out(150) => 
        \data_f0_out[150]\, data_f0_out(149) => 
        \data_f0_out[149]\, data_f0_out(148) => 
        \data_f0_out[148]\, data_f0_out(147) => 
        \data_f0_out[147]\, data_f0_out(146) => 
        \data_f0_out[146]\, data_f0_out(145) => 
        \data_f0_out[145]\, data_f0_out(144) => 
        \data_f0_out[144]\, data_f0_out(143) => 
        \data_f0_out[143]\, data_f0_out(142) => 
        \data_f0_out[142]\, data_f0_out(141) => 
        \data_f0_out[141]\, data_f0_out(140) => 
        \data_f0_out[140]\, data_f0_out(139) => 
        \data_f0_out[139]\, data_f0_out(138) => 
        \data_f0_out[138]\, data_f0_out(137) => 
        \data_f0_out[137]\, data_f0_out(136) => 
        \data_f0_out[136]\, data_f0_out(135) => 
        \data_f0_out[135]\, data_f0_out(134) => 
        \data_f0_out[134]\, data_f0_out(133) => 
        \data_f0_out[133]\, data_f0_out(132) => 
        \data_f0_out[132]\, data_f0_out(131) => 
        \data_f0_out[131]\, data_f0_out(130) => 
        \data_f0_out[130]\, data_f0_out(129) => 
        \data_f0_out[129]\, data_f0_out(128) => 
        \data_f0_out[128]\, data_f0_out(127) => 
        \data_f0_out[127]\, data_f0_out(126) => 
        \data_f0_out[126]\, data_f0_out(125) => 
        \data_f0_out[125]\, data_f0_out(124) => 
        \data_f0_out[124]\, data_f0_out(123) => 
        \data_f0_out[123]\, data_f0_out(122) => 
        \data_f0_out[122]\, data_f0_out(121) => 
        \data_f0_out[121]\, data_f0_out(120) => 
        \data_f0_out[120]\, data_f0_out(119) => 
        \data_f0_out[119]\, data_f0_out(118) => 
        \data_f0_out[118]\, data_f0_out(117) => 
        \data_f0_out[117]\, data_f0_out(116) => 
        \data_f0_out[116]\, data_f0_out(115) => 
        \data_f0_out[115]\, data_f0_out(114) => 
        \data_f0_out[114]\, data_f0_out(113) => 
        \data_f0_out[113]\, data_f0_out(112) => 
        \data_f0_out[112]\, data_f0_out(111) => 
        \data_f0_out[111]\, data_f0_out(110) => 
        \data_f0_out[110]\, data_f0_out(109) => 
        \data_f0_out[109]\, data_f0_out(108) => 
        \data_f0_out[108]\, data_f0_out(107) => 
        \data_f0_out[107]\, data_f0_out(106) => 
        \data_f0_out[106]\, data_f0_out(105) => 
        \data_f0_out[105]\, data_f0_out(104) => 
        \data_f0_out[104]\, data_f0_out(103) => 
        \data_f0_out[103]\, data_f0_out(102) => 
        \data_f0_out[102]\, data_f0_out(101) => 
        \data_f0_out[101]\, data_f0_out(100) => 
        \data_f0_out[100]\, data_f0_out(99) => \data_f0_out[99]\, 
        data_f0_out(98) => \data_f0_out[98]\, data_f0_out(97) => 
        \data_f0_out[97]\, data_f0_out(96) => \data_f0_out[96]\, 
        data_f0_out(95) => \data_f0_out[95]\, data_f0_out(94) => 
        \data_f0_out[94]\, data_f0_out(93) => \data_f0_out[93]\, 
        data_f0_out(92) => \data_f0_out[92]\, data_f0_out(91) => 
        \data_f0_out[91]\, data_f0_out(90) => \data_f0_out[90]\, 
        data_f0_out(89) => \data_f0_out[89]\, data_f0_out(88) => 
        \data_f0_out[88]\, data_f0_out(87) => \data_f0_out[87]\, 
        data_f0_out(86) => \data_f0_out[86]\, data_f0_out(85) => 
        \data_f0_out[85]\, data_f0_out(84) => \data_f0_out[84]\, 
        data_f0_out(83) => \data_f0_out[83]\, data_f0_out(82) => 
        \data_f0_out[82]\, data_f0_out(81) => \data_f0_out[81]\, 
        data_f0_out(80) => \data_f0_out[80]\, data_f0_out(79) => 
        \data_f0_out[79]\, data_f0_out(78) => \data_f0_out[78]\, 
        data_f0_out(77) => \data_f0_out[77]\, data_f0_out(76) => 
        \data_f0_out[76]\, data_f0_out(75) => \data_f0_out[75]\, 
        data_f0_out(74) => \data_f0_out[74]\, data_f0_out(73) => 
        \data_f0_out[73]\, data_f0_out(72) => \data_f0_out[72]\, 
        data_f0_out(71) => \data_f0_out[71]\, data_f0_out(70) => 
        \data_f0_out[70]\, data_f0_out(69) => \data_f0_out[69]\, 
        data_f0_out(68) => \data_f0_out[68]\, data_f0_out(67) => 
        \data_f0_out[67]\, data_f0_out(66) => \data_f0_out[66]\, 
        data_f0_out(65) => \data_f0_out[65]\, data_f0_out(64) => 
        \data_f0_out[64]\, nb_snapshot_param(10) => 
        nb_snapshot_param(10), nb_snapshot_param(9) => 
        nb_snapshot_param(9), nb_snapshot_param(8) => 
        nb_snapshot_param(8), nb_snapshot_param(7) => 
        nb_snapshot_param(7), nb_snapshot_param(6) => 
        nb_snapshot_param(6), nb_snapshot_param(5) => 
        nb_snapshot_param(5), nb_snapshot_param(4) => 
        nb_snapshot_param(4), nb_snapshot_param(3) => 
        nb_snapshot_param(3), nb_snapshot_param(2) => 
        nb_snapshot_param(2), nb_snapshot_param(1) => 
        nb_snapshot_param(1), nb_snapshot_param(0) => 
        nb_snapshot_param(0), sample_f0_37 => sample_f0_37, 
        sample_f0_5 => sample_f0_5, sample_f0_38 => sample_f0_38, 
        sample_f0_6 => sample_f0_6, sample_f0_39 => sample_f0_39, 
        sample_f0_7 => sample_f0_7, sample_f0_40 => sample_f0_40, 
        sample_f0_8 => sample_f0_8, sample_f0_41 => sample_f0_41, 
        sample_f0_9 => sample_f0_9, sample_f0_42 => sample_f0_42, 
        sample_f0_10 => sample_f0_10, sample_f0_43 => 
        sample_f0_43, sample_f0_11 => sample_f0_11, sample_f0_61
         => sample_f0_61, sample_f0_62 => sample_f0_62, 
        sample_f0_63 => sample_f0_63, sample_f0_32 => 
        sample_f0_32, sample_f0_0 => sample_f0_0, sample_f0_33
         => sample_f0_33, sample_f0_1 => sample_f0_1, 
        sample_f0_34 => sample_f0_34, sample_f0_2 => sample_f0_2, 
        sample_f0_35 => sample_f0_35, sample_f0_3 => sample_f0_3, 
        sample_f0_36 => sample_f0_36, sample_f0_4 => sample_f0_4, 
        sample_f0_48 => sample_f0_48, sample_f0_49 => 
        sample_f0_49, sample_f0_50 => sample_f0_50, sample_f0_51
         => sample_f0_51, sample_f0_52 => sample_f0_52, 
        sample_f0_53 => sample_f0_53, sample_f0_54 => 
        sample_f0_54, sample_f0_55 => sample_f0_55, sample_f0_56
         => sample_f0_56, sample_f0_57 => sample_f0_57, 
        sample_f0_58 => sample_f0_58, sample_f0_59 => 
        sample_f0_59, sample_f0_60 => sample_f0_60, sample_f0_44
         => sample_f0_44, sample_f0_12 => sample_f0_12, 
        sample_f0_45 => sample_f0_45, sample_f0_13 => 
        sample_f0_13, sample_f0_46 => sample_f0_46, sample_f0_14
         => sample_f0_14, sample_f0_47 => sample_f0_47, 
        sample_f0_15 => sample_f0_15, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, data_f0_out_valid => data_f0_out_valid, 
        enable_f0 => enable_f0, data_shaping_R0 => 
        data_shaping_R0, data_shaping_R0_0 => data_shaping_R0_0, 
        start_snapshot_f0 => start_snapshot_f0, sample_f0_val_0
         => sample_f0_val_0, burst_f0 => burst_f0);
    
    un7_nb_snapshot_param_more_one_I_31 : XOR2
      port map(A => N_29, B => nb_snapshot_param(6), Y => I_31_5);
    
    lpp_waveform_snapshot_f2 : 
        lpp_waveform_snapshot_160_12_lpp_waveform_snapshot_f1_1
      port map(sample_f2_wdata(95) => sample_f2_wdata(95), 
        sample_f2_wdata(94) => sample_f2_wdata(94), 
        sample_f2_wdata(93) => sample_f2_wdata(93), 
        sample_f2_wdata(92) => sample_f2_wdata(92), 
        sample_f2_wdata(91) => sample_f2_wdata(91), 
        sample_f2_wdata(90) => sample_f2_wdata(90), 
        sample_f2_wdata(89) => sample_f2_wdata(89), 
        sample_f2_wdata(88) => sample_f2_wdata(88), 
        sample_f2_wdata(87) => sample_f2_wdata(87), 
        sample_f2_wdata(86) => sample_f2_wdata(86), 
        sample_f2_wdata(85) => sample_f2_wdata(85), 
        sample_f2_wdata(84) => sample_f2_wdata(84), 
        sample_f2_wdata(83) => sample_f2_wdata(83), 
        sample_f2_wdata(82) => sample_f2_wdata(82), 
        sample_f2_wdata(81) => sample_f2_wdata(81), 
        sample_f2_wdata(80) => sample_f2_wdata(80), 
        sample_f2_wdata(79) => sample_f2_wdata(79), 
        sample_f2_wdata(78) => sample_f2_wdata(78), 
        sample_f2_wdata(77) => sample_f2_wdata(77), 
        sample_f2_wdata(76) => sample_f2_wdata(76), 
        sample_f2_wdata(75) => sample_f2_wdata(75), 
        sample_f2_wdata(74) => sample_f2_wdata(74), 
        sample_f2_wdata(73) => sample_f2_wdata(73), 
        sample_f2_wdata(72) => sample_f2_wdata(72), 
        sample_f2_wdata(71) => sample_f2_wdata(71), 
        sample_f2_wdata(70) => sample_f2_wdata(70), 
        sample_f2_wdata(69) => sample_f2_wdata(69), 
        sample_f2_wdata(68) => sample_f2_wdata(68), 
        sample_f2_wdata(67) => sample_f2_wdata(67), 
        sample_f2_wdata(66) => sample_f2_wdata(66), 
        sample_f2_wdata(65) => sample_f2_wdata(65), 
        sample_f2_wdata(64) => sample_f2_wdata(64), 
        sample_f2_wdata(63) => sample_f2_wdata(63), 
        sample_f2_wdata(62) => sample_f2_wdata(62), 
        sample_f2_wdata(61) => sample_f2_wdata(61), 
        sample_f2_wdata(60) => sample_f2_wdata(60), 
        sample_f2_wdata(59) => sample_f2_wdata(59), 
        sample_f2_wdata(58) => sample_f2_wdata(58), 
        sample_f2_wdata(57) => sample_f2_wdata(57), 
        sample_f2_wdata(56) => sample_f2_wdata(56), 
        sample_f2_wdata(55) => sample_f2_wdata(55), 
        sample_f2_wdata(54) => sample_f2_wdata(54), 
        sample_f2_wdata(53) => sample_f2_wdata(53), 
        sample_f2_wdata(52) => sample_f2_wdata(52), 
        sample_f2_wdata(51) => sample_f2_wdata(51), 
        sample_f2_wdata(50) => sample_f2_wdata(50), 
        sample_f2_wdata(49) => sample_f2_wdata(49), 
        sample_f2_wdata(48) => sample_f2_wdata(48), 
        sample_f2_wdata(47) => sample_f2_wdata(47), 
        sample_f2_wdata(46) => sample_f2_wdata(46), 
        sample_f2_wdata(45) => sample_f2_wdata(45), 
        sample_f2_wdata(44) => sample_f2_wdata(44), 
        sample_f2_wdata(43) => sample_f2_wdata(43), 
        sample_f2_wdata(42) => sample_f2_wdata(42), 
        sample_f2_wdata(41) => sample_f2_wdata(41), 
        sample_f2_wdata(40) => sample_f2_wdata(40), 
        sample_f2_wdata(39) => sample_f2_wdata(39), 
        sample_f2_wdata(38) => sample_f2_wdata(38), 
        sample_f2_wdata(37) => sample_f2_wdata(37), 
        sample_f2_wdata(36) => sample_f2_wdata(36), 
        sample_f2_wdata(35) => sample_f2_wdata(35), 
        sample_f2_wdata(34) => sample_f2_wdata(34), 
        sample_f2_wdata(33) => sample_f2_wdata(33), 
        sample_f2_wdata(32) => sample_f2_wdata(32), 
        sample_f2_wdata(31) => sample_f2_wdata(31), 
        sample_f2_wdata(30) => sample_f2_wdata(30), 
        sample_f2_wdata(29) => sample_f2_wdata(29), 
        sample_f2_wdata(28) => sample_f2_wdata(28), 
        sample_f2_wdata(27) => sample_f2_wdata(27), 
        sample_f2_wdata(26) => sample_f2_wdata(26), 
        sample_f2_wdata(25) => sample_f2_wdata(25), 
        sample_f2_wdata(24) => sample_f2_wdata(24), 
        sample_f2_wdata(23) => sample_f2_wdata(23), 
        sample_f2_wdata(22) => sample_f2_wdata(22), 
        sample_f2_wdata(21) => sample_f2_wdata(21), 
        sample_f2_wdata(20) => sample_f2_wdata(20), 
        sample_f2_wdata(19) => sample_f2_wdata(19), 
        sample_f2_wdata(18) => sample_f2_wdata(18), 
        sample_f2_wdata(17) => sample_f2_wdata(17), 
        sample_f2_wdata(16) => sample_f2_wdata(16), 
        sample_f2_wdata(15) => sample_f2_wdata(15), 
        sample_f2_wdata(14) => sample_f2_wdata(14), 
        sample_f2_wdata(13) => sample_f2_wdata(13), 
        sample_f2_wdata(12) => sample_f2_wdata(12), 
        sample_f2_wdata(11) => sample_f2_wdata(11), 
        sample_f2_wdata(10) => sample_f2_wdata(10), 
        sample_f2_wdata(9) => sample_f2_wdata(9), 
        sample_f2_wdata(8) => sample_f2_wdata(8), 
        sample_f2_wdata(7) => sample_f2_wdata(7), 
        sample_f2_wdata(6) => sample_f2_wdata(6), 
        sample_f2_wdata(5) => sample_f2_wdata(5), 
        sample_f2_wdata(4) => sample_f2_wdata(4), 
        sample_f2_wdata(3) => sample_f2_wdata(3), 
        sample_f2_wdata(2) => sample_f2_wdata(2), 
        sample_f2_wdata(1) => sample_f2_wdata(1), 
        sample_f2_wdata(0) => sample_f2_wdata(0), 
        data_f2_out(159) => \data_f2_out[159]\, data_f2_out(158)
         => \data_f2_out[158]\, data_f2_out(157) => 
        \data_f2_out[157]\, data_f2_out(156) => 
        \data_f2_out[156]\, data_f2_out(155) => 
        \data_f2_out[155]\, data_f2_out(154) => 
        \data_f2_out[154]\, data_f2_out(153) => 
        \data_f2_out[153]\, data_f2_out(152) => 
        \data_f2_out[152]\, data_f2_out(151) => 
        \data_f2_out[151]\, data_f2_out(150) => 
        \data_f2_out[150]\, data_f2_out(149) => 
        \data_f2_out[149]\, data_f2_out(148) => 
        \data_f2_out[148]\, data_f2_out(147) => 
        \data_f2_out[147]\, data_f2_out(146) => 
        \data_f2_out[146]\, data_f2_out(145) => 
        \data_f2_out[145]\, data_f2_out(144) => 
        \data_f2_out[144]\, data_f2_out(143) => 
        \data_f2_out[143]\, data_f2_out(142) => 
        \data_f2_out[142]\, data_f2_out(141) => 
        \data_f2_out[141]\, data_f2_out(140) => 
        \data_f2_out[140]\, data_f2_out(139) => 
        \data_f2_out[139]\, data_f2_out(138) => 
        \data_f2_out[138]\, data_f2_out(137) => 
        \data_f2_out[137]\, data_f2_out(136) => 
        \data_f2_out[136]\, data_f2_out(135) => 
        \data_f2_out[135]\, data_f2_out(134) => 
        \data_f2_out[134]\, data_f2_out(133) => 
        \data_f2_out[133]\, data_f2_out(132) => 
        \data_f2_out[132]\, data_f2_out(131) => 
        \data_f2_out[131]\, data_f2_out(130) => 
        \data_f2_out[130]\, data_f2_out(129) => 
        \data_f2_out[129]\, data_f2_out(128) => 
        \data_f2_out[128]\, data_f2_out(127) => 
        \data_f2_out[127]\, data_f2_out(126) => 
        \data_f2_out[126]\, data_f2_out(125) => 
        \data_f2_out[125]\, data_f2_out(124) => 
        \data_f2_out[124]\, data_f2_out(123) => 
        \data_f2_out[123]\, data_f2_out(122) => 
        \data_f2_out[122]\, data_f2_out(121) => 
        \data_f2_out[121]\, data_f2_out(120) => 
        \data_f2_out[120]\, data_f2_out(119) => 
        \data_f2_out[119]\, data_f2_out(118) => 
        \data_f2_out[118]\, data_f2_out(117) => 
        \data_f2_out[117]\, data_f2_out(116) => 
        \data_f2_out[116]\, data_f2_out(115) => 
        \data_f2_out[115]\, data_f2_out(114) => 
        \data_f2_out[114]\, data_f2_out(113) => 
        \data_f2_out[113]\, data_f2_out(112) => 
        \data_f2_out[112]\, data_f2_out(111) => 
        \data_f2_out[111]\, data_f2_out(110) => 
        \data_f2_out[110]\, data_f2_out(109) => 
        \data_f2_out[109]\, data_f2_out(108) => 
        \data_f2_out[108]\, data_f2_out(107) => 
        \data_f2_out[107]\, data_f2_out(106) => 
        \data_f2_out[106]\, data_f2_out(105) => 
        \data_f2_out[105]\, data_f2_out(104) => 
        \data_f2_out[104]\, data_f2_out(103) => 
        \data_f2_out[103]\, data_f2_out(102) => 
        \data_f2_out[102]\, data_f2_out(101) => 
        \data_f2_out[101]\, data_f2_out(100) => 
        \data_f2_out[100]\, data_f2_out(99) => \data_f2_out[99]\, 
        data_f2_out(98) => \data_f2_out[98]\, data_f2_out(97) => 
        \data_f2_out[97]\, data_f2_out(96) => \data_f2_out[96]\, 
        data_f2_out(95) => \data_f2_out[95]\, data_f2_out(94) => 
        \data_f2_out[94]\, data_f2_out(93) => \data_f2_out[93]\, 
        data_f2_out(92) => \data_f2_out[92]\, data_f2_out(91) => 
        \data_f2_out[91]\, data_f2_out(90) => \data_f2_out[90]\, 
        data_f2_out(89) => \data_f2_out[89]\, data_f2_out(88) => 
        \data_f2_out[88]\, data_f2_out(87) => \data_f2_out[87]\, 
        data_f2_out(86) => \data_f2_out[86]\, data_f2_out(85) => 
        \data_f2_out[85]\, data_f2_out(84) => \data_f2_out[84]\, 
        data_f2_out(83) => \data_f2_out[83]\, data_f2_out(82) => 
        \data_f2_out[82]\, data_f2_out(81) => \data_f2_out[81]\, 
        data_f2_out(80) => \data_f2_out[80]\, data_f2_out(79) => 
        \data_f2_out[79]\, data_f2_out(78) => \data_f2_out[78]\, 
        data_f2_out(77) => \data_f2_out[77]\, data_f2_out(76) => 
        \data_f2_out[76]\, data_f2_out(75) => \data_f2_out[75]\, 
        data_f2_out(74) => \data_f2_out[74]\, data_f2_out(73) => 
        \data_f2_out[73]\, data_f2_out(72) => \data_f2_out[72]\, 
        data_f2_out(71) => \data_f2_out[71]\, data_f2_out(70) => 
        \data_f2_out[70]\, data_f2_out(69) => \data_f2_out[69]\, 
        data_f2_out(68) => \data_f2_out[68]\, data_f2_out(67) => 
        \data_f2_out[67]\, data_f2_out(66) => \data_f2_out[66]\, 
        data_f2_out(65) => \data_f2_out[65]\, data_f2_out(64) => 
        \data_f2_out[64]\, nb_snapshot_param(0) => 
        nb_snapshot_param(0), HRESETn_c => HRESETn_c, HCLK_c => 
        HCLK_c, data_f2_out_valid => data_f2_out_valid, I_13_20
         => I_13_20, I_9_20 => I_9_20, I_5_20 => I_5_20, I_38_4
         => I_38_4, I_31_5 => I_31_5, N_4 => N_4, I_45_4 => 
        I_45_4, I_56_4 => I_56_4, I_52_4 => I_52_4, I_24_4 => 
        I_24_4, I_20_12 => I_20_12, enable_f2 => enable_f2, 
        burst_f2 => burst_f2, start_snapshot_f2 => 
        start_snapshot_f2, sample_f2_val => sample_f2_val);
    
    un7_nb_snapshot_param_more_one_I_12 : AND3
      port map(A => nb_snapshot_param(0), B => 
        nb_snapshot_param(1), C => nb_snapshot_param(2), Y => 
        N_42);
    
    un7_nb_snapshot_param_more_one_I_5 : XOR2
      port map(A => nb_snapshot_param(0), B => 
        nb_snapshot_param(1), Y => I_5_20);
    
    un7_nb_snapshot_param_more_one_I_51 : NOR2B
      port map(A => nb_snapshot_param(8), B => \DWACT_FINC_E[4]\, 
        Y => N_14);
    
    pp_waveform_dma_1 : lpp_waveform_dma
      port map(addr_data_f0(31) => addr_data_f0(31), 
        addr_data_f0(30) => addr_data_f0(30), addr_data_f0(29)
         => addr_data_f0(29), addr_data_f0(28) => 
        addr_data_f0(28), addr_data_f0(27) => addr_data_f0(27), 
        addr_data_f0(26) => addr_data_f0(26), addr_data_f0(25)
         => addr_data_f0(25), addr_data_f0(24) => 
        addr_data_f0(24), addr_data_f0(23) => addr_data_f0(23), 
        addr_data_f0(22) => addr_data_f0(22), addr_data_f0(21)
         => addr_data_f0(21), addr_data_f0(20) => 
        addr_data_f0(20), addr_data_f0(19) => addr_data_f0(19), 
        addr_data_f0(18) => addr_data_f0(18), addr_data_f0(17)
         => addr_data_f0(17), addr_data_f0(16) => 
        addr_data_f0(16), addr_data_f0(15) => addr_data_f0(15), 
        addr_data_f0(14) => addr_data_f0(14), addr_data_f0(13)
         => addr_data_f0(13), addr_data_f0(12) => 
        addr_data_f0(12), addr_data_f0(11) => addr_data_f0(11), 
        addr_data_f0(10) => addr_data_f0(10), addr_data_f0(9) => 
        addr_data_f0(9), addr_data_f0(8) => addr_data_f0(8), 
        addr_data_f0(7) => addr_data_f0(7), addr_data_f0(6) => 
        addr_data_f0(6), addr_data_f0(5) => addr_data_f0(5), 
        addr_data_f0(4) => addr_data_f0(4), addr_data_f0(3) => 
        addr_data_f0(3), addr_data_f0(2) => addr_data_f0(2), 
        addr_data_f0(1) => addr_data_f0(1), addr_data_f0(0) => 
        addr_data_f0(0), addr_data_f1(31) => addr_data_f1(31), 
        addr_data_f1(30) => addr_data_f1(30), addr_data_f1(29)
         => addr_data_f1(29), addr_data_f1(28) => 
        addr_data_f1(28), addr_data_f1(27) => addr_data_f1(27), 
        addr_data_f1(26) => addr_data_f1(26), addr_data_f1(25)
         => addr_data_f1(25), addr_data_f1(24) => 
        addr_data_f1(24), addr_data_f1(23) => addr_data_f1(23), 
        addr_data_f1(22) => addr_data_f1(22), addr_data_f1(21)
         => addr_data_f1(21), addr_data_f1(20) => 
        addr_data_f1(20), addr_data_f1(19) => addr_data_f1(19), 
        addr_data_f1(18) => addr_data_f1(18), addr_data_f1(17)
         => addr_data_f1(17), addr_data_f1(16) => 
        addr_data_f1(16), addr_data_f1(15) => addr_data_f1(15), 
        addr_data_f1(14) => addr_data_f1(14), addr_data_f1(13)
         => addr_data_f1(13), addr_data_f1(12) => 
        addr_data_f1(12), addr_data_f1(11) => addr_data_f1(11), 
        addr_data_f1(10) => addr_data_f1(10), addr_data_f1(9) => 
        addr_data_f1(9), addr_data_f1(8) => addr_data_f1(8), 
        addr_data_f1(7) => addr_data_f1(7), addr_data_f1(6) => 
        addr_data_f1(6), addr_data_f1(5) => addr_data_f1(5), 
        addr_data_f1(4) => addr_data_f1(4), addr_data_f1(3) => 
        addr_data_f1(3), addr_data_f1(2) => addr_data_f1(2), 
        addr_data_f1(1) => addr_data_f1(1), addr_data_f1(0) => 
        addr_data_f1(0), addr_data_f2(31) => addr_data_f2(31), 
        addr_data_f2(30) => addr_data_f2(30), addr_data_f2(29)
         => addr_data_f2(29), addr_data_f2(28) => 
        addr_data_f2(28), addr_data_f2(27) => addr_data_f2(27), 
        addr_data_f2(26) => addr_data_f2(26), addr_data_f2(25)
         => addr_data_f2(25), addr_data_f2(24) => 
        addr_data_f2(24), addr_data_f2(23) => addr_data_f2(23), 
        addr_data_f2(22) => addr_data_f2(22), addr_data_f2(21)
         => addr_data_f2(21), addr_data_f2(20) => 
        addr_data_f2(20), addr_data_f2(19) => addr_data_f2(19), 
        addr_data_f2(18) => addr_data_f2(18), addr_data_f2(17)
         => addr_data_f2(17), addr_data_f2(16) => 
        addr_data_f2(16), addr_data_f2(15) => addr_data_f2(15), 
        addr_data_f2(14) => addr_data_f2(14), addr_data_f2(13)
         => addr_data_f2(13), addr_data_f2(12) => 
        addr_data_f2(12), addr_data_f2(11) => addr_data_f2(11), 
        addr_data_f2(10) => addr_data_f2(10), addr_data_f2(9) => 
        addr_data_f2(9), addr_data_f2(8) => addr_data_f2(8), 
        addr_data_f2(7) => addr_data_f2(7), addr_data_f2(6) => 
        addr_data_f2(6), addr_data_f2(5) => addr_data_f2(5), 
        addr_data_f2(4) => addr_data_f2(4), addr_data_f2(3) => 
        addr_data_f2(3), addr_data_f2(2) => addr_data_f2(2), 
        addr_data_f2(1) => addr_data_f2(1), addr_data_f2(0) => 
        addr_data_f2(0), addr_data_f3(31) => addr_data_f3(31), 
        addr_data_f3(30) => addr_data_f3(30), addr_data_f3(29)
         => addr_data_f3(29), addr_data_f3(28) => 
        addr_data_f3(28), addr_data_f3(27) => addr_data_f3(27), 
        addr_data_f3(26) => addr_data_f3(26), addr_data_f3(25)
         => addr_data_f3(25), addr_data_f3(24) => 
        addr_data_f3(24), addr_data_f3(23) => addr_data_f3(23), 
        addr_data_f3(22) => addr_data_f3(22), addr_data_f3(21)
         => addr_data_f3(21), addr_data_f3(20) => 
        addr_data_f3(20), addr_data_f3(19) => addr_data_f3(19), 
        addr_data_f3(18) => addr_data_f3(18), addr_data_f3(17)
         => addr_data_f3(17), addr_data_f3(16) => 
        addr_data_f3(16), addr_data_f3(15) => addr_data_f3(15), 
        addr_data_f3(14) => addr_data_f3(14), addr_data_f3(13)
         => addr_data_f3(13), addr_data_f3(12) => 
        addr_data_f3(12), addr_data_f3(11) => addr_data_f3(11), 
        addr_data_f3(10) => addr_data_f3(10), addr_data_f3(9) => 
        addr_data_f3(9), addr_data_f3(8) => addr_data_f3(8), 
        addr_data_f3(7) => addr_data_f3(7), addr_data_f3(6) => 
        addr_data_f3(6), addr_data_f3(5) => addr_data_f3(5), 
        addr_data_f3(4) => addr_data_f3(4), addr_data_f3(3) => 
        addr_data_f3(3), addr_data_f3(2) => addr_data_f3(2), 
        addr_data_f3(1) => addr_data_f3(1), addr_data_f3(0) => 
        addr_data_f3(0), status_full(3) => status_full(3), 
        status_full(2) => status_full(2), status_full(1) => 
        status_full(1), status_full(0) => status_full(0), 
        status_full_err(3) => status_full_err(3), 
        status_full_err(2) => status_full_err(2), 
        status_full_err(1) => status_full_err(1), 
        status_full_err(0) => status_full_err(0), 
        nb_burst_available(10) => nb_burst_available(10), 
        nb_burst_available(9) => nb_burst_available(9), 
        nb_burst_available(8) => nb_burst_available(8), 
        nb_burst_available(7) => nb_burst_available(7), 
        nb_burst_available(6) => nb_burst_available(6), 
        nb_burst_available(5) => nb_burst_available(5), 
        nb_burst_available(4) => nb_burst_available(4), 
        nb_burst_available(3) => nb_burst_available(3), 
        nb_burst_available(2) => nb_burst_available(2), 
        nb_burst_available(1) => nb_burst_available(1), 
        nb_burst_available(0) => nb_burst_available(0), 
        haddr_c(31) => haddr_c(31), haddr_c(30) => haddr_c(30), 
        haddr_c(29) => haddr_c(29), haddr_c(28) => haddr_c(28), 
        haddr_c(27) => haddr_c(27), haddr_c(26) => haddr_c(26), 
        haddr_c(25) => haddr_c(25), haddr_c(24) => haddr_c(24), 
        haddr_c(23) => haddr_c(23), haddr_c(22) => haddr_c(22), 
        haddr_c(21) => haddr_c(21), haddr_c(20) => haddr_c(20), 
        haddr_c(19) => haddr_c(19), haddr_c(18) => haddr_c(18), 
        haddr_c(17) => haddr_c(17), haddr_c(16) => haddr_c(16), 
        haddr_c(15) => haddr_c(15), haddr_c(14) => haddr_c(14), 
        haddr_c(13) => haddr_c(13), haddr_c(12) => haddr_c(12), 
        haddr_c(11) => haddr_c(11), haddr_c(10) => haddr_c(10), 
        haddr_c(9) => haddr_c(9), haddr_c(8) => haddr_c(8), 
        haddr_c(7) => haddr_c(7), haddr_c(6) => haddr_c(6), 
        haddr_c(5) => haddr_c(5), haddr_c(4) => haddr_c(4), 
        haddr_c(3) => haddr_c(3), haddr_c(2) => haddr_c(2), 
        haddr_c(1) => haddr_c(1), haddr_c(0) => haddr_c(0), 
        AHB_Master_In_c_3 => AHB_Master_In_c_3, AHB_Master_In_c_0
         => AHB_Master_In_c_0, AHB_Master_In_c_4 => 
        AHB_Master_In_c_4, AHB_Master_In_c_5 => AHB_Master_In_c_5, 
        hsize_c(1) => hsize_c(1), hsize_c(0) => hsize_c(0), 
        htrans_c(1) => htrans_c(1), htrans_c(0) => htrans_c(0), 
        hburst_c(2) => hburst_c(2), hburst_c(1) => hburst_c(1), 
        hburst_c(0) => hburst_c(0), status_full_ack(3) => 
        status_full_ack(3), status_full_ack(2) => 
        status_full_ack(2), status_full_ack(1) => 
        status_full_ack(1), status_full_ack(0) => 
        status_full_ack(0), ready_i_0(3) => \ready_i_0[3]\, 
        ready_i_0(2) => \ready_i_0[2]\, ready_i_0(1) => 
        \ready_i_0[1]\, ready_i_0(0) => \ready_i_0[0]\, 
        data_ren(3) => \data_ren[3]\, data_ren(2) => 
        \data_ren[2]\, data_ren(1) => \data_ren[1]\, data_ren(0)
         => \data_ren[0]\, time_ren(3) => \time_ren[3]\, 
        time_ren(2) => \time_ren[2]\, time_ren(1) => 
        \time_ren[1]\, time_ren(0) => \time_ren[0]\, time_ren_1z
         => time_ren, data_ren_1z => data_ren, N_43 => N_43, 
        IdlePhase_RNI03G71 => IdlePhase_RNI03G71, hwrite_c => 
        hwrite_c, un20_time_write => un20_time_write, 
        un13_time_write => un13_time_write, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c);
    
    lpp_waveform_fifo_arbiter_1 : lpp_waveform_fifo_arbiter
      port map(wdata(31) => \wdata[31]\, wdata(30) => \wdata[30]\, 
        wdata(29) => \wdata[29]\, wdata(28) => \wdata[28]\, 
        wdata(27) => \wdata[27]\, wdata(26) => \wdata[26]\, 
        wdata(25) => \wdata[25]\, wdata(24) => \wdata[24]\, 
        wdata(23) => \wdata[23]\, wdata(22) => \wdata[22]\, 
        wdata(21) => \wdata[21]\, wdata(20) => \wdata[20]\, 
        wdata(19) => \wdata[19]\, wdata(18) => \wdata[18]\, 
        wdata(17) => \wdata[17]\, wdata(16) => \wdata[16]\, 
        wdata(15) => \wdata[15]\, wdata(14) => \wdata[14]\, 
        wdata(13) => \wdata[13]\, wdata(12) => \wdata[12]\, 
        wdata(11) => \wdata[11]\, wdata(10) => \wdata[10]\, 
        wdata(9) => \wdata[9]\, wdata(8) => \wdata[8]\, wdata(7)
         => \wdata[7]\, wdata(6) => \wdata[6]\, wdata(5) => 
        \wdata[5]\, wdata(4) => \wdata[4]\, wdata(3) => 
        \wdata[3]\, wdata(2) => \wdata[2]\, wdata(1) => 
        \wdata[1]\, wdata(0) => \wdata[0]\, data_wen(3) => 
        \data_wen[3]\, data_wen(2) => \data_wen[2]\, data_wen(1)
         => \data_wen[1]\, data_wen(0) => \data_wen[0]\, 
        valid_ack(3) => \valid_ack[3]\, valid_ack(2) => 
        \valid_ack[2]\, valid_ack(1) => \valid_ack[1]\, 
        valid_ack(0) => \valid_ack[0]\, time_wen(3) => 
        \time_wen[3]\, time_wen(2) => \time_wen[2]\, time_wen(1)
         => \time_wen[1]\, time_wen(0) => \time_wen[0]\, 
        data_f3_out(159) => \data_f3_out[159]\, data_f3_out(158)
         => \data_f3_out[158]\, data_f3_out(157) => 
        \data_f3_out[157]\, data_f3_out(156) => 
        \data_f3_out[156]\, data_f3_out(155) => 
        \data_f3_out[155]\, data_f3_out(154) => 
        \data_f3_out[154]\, data_f3_out(153) => 
        \data_f3_out[153]\, data_f3_out(152) => 
        \data_f3_out[152]\, data_f3_out(151) => 
        \data_f3_out[151]\, data_f3_out(150) => 
        \data_f3_out[150]\, data_f3_out(149) => 
        \data_f3_out[149]\, data_f3_out(148) => 
        \data_f3_out[148]\, data_f3_out(147) => 
        \data_f3_out[147]\, data_f3_out(146) => 
        \data_f3_out[146]\, data_f3_out(145) => 
        \data_f3_out[145]\, data_f3_out(144) => 
        \data_f3_out[144]\, data_f3_out(143) => 
        \data_f3_out[143]\, data_f3_out(142) => 
        \data_f3_out[142]\, data_f3_out(141) => 
        \data_f3_out[141]\, data_f3_out(140) => 
        \data_f3_out[140]\, data_f3_out(139) => 
        \data_f3_out[139]\, data_f3_out(138) => 
        \data_f3_out[138]\, data_f3_out(137) => 
        \data_f3_out[137]\, data_f3_out(136) => 
        \data_f3_out[136]\, data_f3_out(135) => 
        \data_f3_out[135]\, data_f3_out(134) => 
        \data_f3_out[134]\, data_f3_out(133) => 
        \data_f3_out[133]\, data_f3_out(132) => 
        \data_f3_out[132]\, data_f3_out(131) => 
        \data_f3_out[131]\, data_f3_out(130) => 
        \data_f3_out[130]\, data_f3_out(129) => 
        \data_f3_out[129]\, data_f3_out(128) => 
        \data_f3_out[128]\, data_f3_out(127) => 
        \data_f3_out[127]\, data_f3_out(126) => 
        \data_f3_out[126]\, data_f3_out(125) => 
        \data_f3_out[125]\, data_f3_out(124) => 
        \data_f3_out[124]\, data_f3_out(123) => 
        \data_f3_out[123]\, data_f3_out(122) => 
        \data_f3_out[122]\, data_f3_out(121) => 
        \data_f3_out[121]\, data_f3_out(120) => 
        \data_f3_out[120]\, data_f3_out(119) => 
        \data_f3_out[119]\, data_f3_out(118) => 
        \data_f3_out[118]\, data_f3_out(117) => 
        \data_f3_out[117]\, data_f3_out(116) => 
        \data_f3_out[116]\, data_f3_out(115) => 
        \data_f3_out[115]\, data_f3_out(114) => 
        \data_f3_out[114]\, data_f3_out(113) => 
        \data_f3_out[113]\, data_f3_out(112) => 
        \data_f3_out[112]\, data_f3_out(111) => 
        \data_f3_out[111]\, data_f3_out(110) => 
        \data_f3_out[110]\, data_f3_out(109) => 
        \data_f3_out[109]\, data_f3_out(108) => 
        \data_f3_out[108]\, data_f3_out(107) => 
        \data_f3_out[107]\, data_f3_out(106) => 
        \data_f3_out[106]\, data_f3_out(105) => 
        \data_f3_out[105]\, data_f3_out(104) => 
        \data_f3_out[104]\, data_f3_out(103) => 
        \data_f3_out[103]\, data_f3_out(102) => 
        \data_f3_out[102]\, data_f3_out(101) => 
        \data_f3_out[101]\, data_f3_out(100) => 
        \data_f3_out[100]\, data_f3_out(99) => \data_f3_out[99]\, 
        data_f3_out(98) => \data_f3_out[98]\, data_f3_out(97) => 
        \data_f3_out[97]\, data_f3_out(96) => \data_f3_out[96]\, 
        data_f3_out(95) => \data_f3_out[95]\, data_f3_out(94) => 
        \data_f3_out[94]\, data_f3_out(93) => \data_f3_out[93]\, 
        data_f3_out(92) => \data_f3_out[92]\, data_f3_out(91) => 
        \data_f3_out[91]\, data_f3_out(90) => \data_f3_out[90]\, 
        data_f3_out(89) => \data_f3_out[89]\, data_f3_out(88) => 
        \data_f3_out[88]\, data_f3_out(87) => \data_f3_out[87]\, 
        data_f3_out(86) => \data_f3_out[86]\, data_f3_out(85) => 
        \data_f3_out[85]\, data_f3_out(84) => \data_f3_out[84]\, 
        data_f3_out(83) => \data_f3_out[83]\, data_f3_out(82) => 
        \data_f3_out[82]\, data_f3_out(81) => \data_f3_out[81]\, 
        data_f3_out(80) => \data_f3_out[80]\, data_f3_out(79) => 
        \data_f3_out[79]\, data_f3_out(78) => \data_f3_out[78]\, 
        data_f3_out(77) => \data_f3_out[77]\, data_f3_out(76) => 
        \data_f3_out[76]\, data_f3_out(75) => \data_f3_out[75]\, 
        data_f3_out(74) => \data_f3_out[74]\, data_f3_out(73) => 
        \data_f3_out[73]\, data_f3_out(72) => \data_f3_out[72]\, 
        data_f3_out(71) => \data_f3_out[71]\, data_f3_out(70) => 
        \data_f3_out[70]\, data_f3_out(69) => \data_f3_out[69]\, 
        data_f3_out(68) => \data_f3_out[68]\, data_f3_out(67) => 
        \data_f3_out[67]\, data_f3_out(66) => \data_f3_out[66]\, 
        data_f3_out(65) => \data_f3_out[65]\, data_f3_out(64) => 
        \data_f3_out[64]\, data_f2_out(159) => \data_f2_out[159]\, 
        data_f2_out(158) => \data_f2_out[158]\, data_f2_out(157)
         => \data_f2_out[157]\, data_f2_out(156) => 
        \data_f2_out[156]\, data_f2_out(155) => 
        \data_f2_out[155]\, data_f2_out(154) => 
        \data_f2_out[154]\, data_f2_out(153) => 
        \data_f2_out[153]\, data_f2_out(152) => 
        \data_f2_out[152]\, data_f2_out(151) => 
        \data_f2_out[151]\, data_f2_out(150) => 
        \data_f2_out[150]\, data_f2_out(149) => 
        \data_f2_out[149]\, data_f2_out(148) => 
        \data_f2_out[148]\, data_f2_out(147) => 
        \data_f2_out[147]\, data_f2_out(146) => 
        \data_f2_out[146]\, data_f2_out(145) => 
        \data_f2_out[145]\, data_f2_out(144) => 
        \data_f2_out[144]\, data_f2_out(143) => 
        \data_f2_out[143]\, data_f2_out(142) => 
        \data_f2_out[142]\, data_f2_out(141) => 
        \data_f2_out[141]\, data_f2_out(140) => 
        \data_f2_out[140]\, data_f2_out(139) => 
        \data_f2_out[139]\, data_f2_out(138) => 
        \data_f2_out[138]\, data_f2_out(137) => 
        \data_f2_out[137]\, data_f2_out(136) => 
        \data_f2_out[136]\, data_f2_out(135) => 
        \data_f2_out[135]\, data_f2_out(134) => 
        \data_f2_out[134]\, data_f2_out(133) => 
        \data_f2_out[133]\, data_f2_out(132) => 
        \data_f2_out[132]\, data_f2_out(131) => 
        \data_f2_out[131]\, data_f2_out(130) => 
        \data_f2_out[130]\, data_f2_out(129) => 
        \data_f2_out[129]\, data_f2_out(128) => 
        \data_f2_out[128]\, data_f2_out(127) => 
        \data_f2_out[127]\, data_f2_out(126) => 
        \data_f2_out[126]\, data_f2_out(125) => 
        \data_f2_out[125]\, data_f2_out(124) => 
        \data_f2_out[124]\, data_f2_out(123) => 
        \data_f2_out[123]\, data_f2_out(122) => 
        \data_f2_out[122]\, data_f2_out(121) => 
        \data_f2_out[121]\, data_f2_out(120) => 
        \data_f2_out[120]\, data_f2_out(119) => 
        \data_f2_out[119]\, data_f2_out(118) => 
        \data_f2_out[118]\, data_f2_out(117) => 
        \data_f2_out[117]\, data_f2_out(116) => 
        \data_f2_out[116]\, data_f2_out(115) => 
        \data_f2_out[115]\, data_f2_out(114) => 
        \data_f2_out[114]\, data_f2_out(113) => 
        \data_f2_out[113]\, data_f2_out(112) => 
        \data_f2_out[112]\, data_f2_out(111) => 
        \data_f2_out[111]\, data_f2_out(110) => 
        \data_f2_out[110]\, data_f2_out(109) => 
        \data_f2_out[109]\, data_f2_out(108) => 
        \data_f2_out[108]\, data_f2_out(107) => 
        \data_f2_out[107]\, data_f2_out(106) => 
        \data_f2_out[106]\, data_f2_out(105) => 
        \data_f2_out[105]\, data_f2_out(104) => 
        \data_f2_out[104]\, data_f2_out(103) => 
        \data_f2_out[103]\, data_f2_out(102) => 
        \data_f2_out[102]\, data_f2_out(101) => 
        \data_f2_out[101]\, data_f2_out(100) => 
        \data_f2_out[100]\, data_f2_out(99) => \data_f2_out[99]\, 
        data_f2_out(98) => \data_f2_out[98]\, data_f2_out(97) => 
        \data_f2_out[97]\, data_f2_out(96) => \data_f2_out[96]\, 
        data_f2_out(95) => \data_f2_out[95]\, data_f2_out(94) => 
        \data_f2_out[94]\, data_f2_out(93) => \data_f2_out[93]\, 
        data_f2_out(92) => \data_f2_out[92]\, data_f2_out(91) => 
        \data_f2_out[91]\, data_f2_out(90) => \data_f2_out[90]\, 
        data_f2_out(89) => \data_f2_out[89]\, data_f2_out(88) => 
        \data_f2_out[88]\, data_f2_out(87) => \data_f2_out[87]\, 
        data_f2_out(86) => \data_f2_out[86]\, data_f2_out(85) => 
        \data_f2_out[85]\, data_f2_out(84) => \data_f2_out[84]\, 
        data_f2_out(83) => \data_f2_out[83]\, data_f2_out(82) => 
        \data_f2_out[82]\, data_f2_out(81) => \data_f2_out[81]\, 
        data_f2_out(80) => \data_f2_out[80]\, data_f2_out(79) => 
        \data_f2_out[79]\, data_f2_out(78) => \data_f2_out[78]\, 
        data_f2_out(77) => \data_f2_out[77]\, data_f2_out(76) => 
        \data_f2_out[76]\, data_f2_out(75) => \data_f2_out[75]\, 
        data_f2_out(74) => \data_f2_out[74]\, data_f2_out(73) => 
        \data_f2_out[73]\, data_f2_out(72) => \data_f2_out[72]\, 
        data_f2_out(71) => \data_f2_out[71]\, data_f2_out(70) => 
        \data_f2_out[70]\, data_f2_out(69) => \data_f2_out[69]\, 
        data_f2_out(68) => \data_f2_out[68]\, data_f2_out(67) => 
        \data_f2_out[67]\, data_f2_out(66) => \data_f2_out[66]\, 
        data_f2_out(65) => \data_f2_out[65]\, data_f2_out(64) => 
        \data_f2_out[64]\, data_f1_out(159) => \data_f1_out[159]\, 
        data_f1_out(158) => \data_f1_out[158]\, data_f1_out(157)
         => \data_f1_out[157]\, data_f1_out(156) => 
        \data_f1_out[156]\, data_f1_out(155) => 
        \data_f1_out[155]\, data_f1_out(154) => 
        \data_f1_out[154]\, data_f1_out(153) => 
        \data_f1_out[153]\, data_f1_out(152) => 
        \data_f1_out[152]\, data_f1_out(151) => 
        \data_f1_out[151]\, data_f1_out(150) => 
        \data_f1_out[150]\, data_f1_out(149) => 
        \data_f1_out[149]\, data_f1_out(148) => 
        \data_f1_out[148]\, data_f1_out(147) => 
        \data_f1_out[147]\, data_f1_out(146) => 
        \data_f1_out[146]\, data_f1_out(145) => 
        \data_f1_out[145]\, data_f1_out(144) => 
        \data_f1_out[144]\, data_f1_out(143) => 
        \data_f1_out[143]\, data_f1_out(142) => 
        \data_f1_out[142]\, data_f1_out(141) => 
        \data_f1_out[141]\, data_f1_out(140) => 
        \data_f1_out[140]\, data_f1_out(139) => 
        \data_f1_out[139]\, data_f1_out(138) => 
        \data_f1_out[138]\, data_f1_out(137) => 
        \data_f1_out[137]\, data_f1_out(136) => 
        \data_f1_out[136]\, data_f1_out(135) => 
        \data_f1_out[135]\, data_f1_out(134) => 
        \data_f1_out[134]\, data_f1_out(133) => 
        \data_f1_out[133]\, data_f1_out(132) => 
        \data_f1_out[132]\, data_f1_out(131) => 
        \data_f1_out[131]\, data_f1_out(130) => 
        \data_f1_out[130]\, data_f1_out(129) => 
        \data_f1_out[129]\, data_f1_out(128) => 
        \data_f1_out[128]\, data_f1_out(127) => 
        \data_f1_out[127]\, data_f1_out(126) => 
        \data_f1_out[126]\, data_f1_out(125) => 
        \data_f1_out[125]\, data_f1_out(124) => 
        \data_f1_out[124]\, data_f1_out(123) => 
        \data_f1_out[123]\, data_f1_out(122) => 
        \data_f1_out[122]\, data_f1_out(121) => 
        \data_f1_out[121]\, data_f1_out(120) => 
        \data_f1_out[120]\, data_f1_out(119) => 
        \data_f1_out[119]\, data_f1_out(118) => 
        \data_f1_out[118]\, data_f1_out(117) => 
        \data_f1_out[117]\, data_f1_out(116) => 
        \data_f1_out[116]\, data_f1_out(115) => 
        \data_f1_out[115]\, data_f1_out(114) => 
        \data_f1_out[114]\, data_f1_out(113) => 
        \data_f1_out[113]\, data_f1_out(112) => 
        \data_f1_out[112]\, data_f1_out(111) => 
        \data_f1_out[111]\, data_f1_out(110) => 
        \data_f1_out[110]\, data_f1_out(109) => 
        \data_f1_out[109]\, data_f1_out(108) => 
        \data_f1_out[108]\, data_f1_out(107) => 
        \data_f1_out[107]\, data_f1_out(106) => 
        \data_f1_out[106]\, data_f1_out(105) => 
        \data_f1_out[105]\, data_f1_out(104) => 
        \data_f1_out[104]\, data_f1_out(103) => 
        \data_f1_out[103]\, data_f1_out(102) => 
        \data_f1_out[102]\, data_f1_out(101) => 
        \data_f1_out[101]\, data_f1_out(100) => 
        \data_f1_out[100]\, data_f1_out(99) => \data_f1_out[99]\, 
        data_f1_out(98) => \data_f1_out[98]\, data_f1_out(97) => 
        \data_f1_out[97]\, data_f1_out(96) => \data_f1_out[96]\, 
        data_f1_out(95) => \data_f1_out[95]\, data_f1_out(94) => 
        \data_f1_out[94]\, data_f1_out(93) => \data_f1_out[93]\, 
        data_f1_out(92) => \data_f1_out[92]\, data_f1_out(91) => 
        \data_f1_out[91]\, data_f1_out(90) => \data_f1_out[90]\, 
        data_f1_out(89) => \data_f1_out[89]\, data_f1_out(88) => 
        \data_f1_out[88]\, data_f1_out(87) => \data_f1_out[87]\, 
        data_f1_out(86) => \data_f1_out[86]\, data_f1_out(85) => 
        \data_f1_out[85]\, data_f1_out(84) => \data_f1_out[84]\, 
        data_f1_out(83) => \data_f1_out[83]\, data_f1_out(82) => 
        \data_f1_out[82]\, data_f1_out(81) => \data_f1_out[81]\, 
        data_f1_out(80) => \data_f1_out[80]\, data_f1_out(79) => 
        \data_f1_out[79]\, data_f1_out(78) => \data_f1_out[78]\, 
        data_f1_out(77) => \data_f1_out[77]\, data_f1_out(76) => 
        \data_f1_out[76]\, data_f1_out(75) => \data_f1_out[75]\, 
        data_f1_out(74) => \data_f1_out[74]\, data_f1_out(73) => 
        \data_f1_out[73]\, data_f1_out(72) => \data_f1_out[72]\, 
        data_f1_out(71) => \data_f1_out[71]\, data_f1_out(70) => 
        \data_f1_out[70]\, data_f1_out(69) => \data_f1_out[69]\, 
        data_f1_out(68) => \data_f1_out[68]\, data_f1_out(67) => 
        \data_f1_out[67]\, data_f1_out(66) => \data_f1_out[66]\, 
        data_f1_out(65) => \data_f1_out[65]\, data_f1_out(64) => 
        \data_f1_out[64]\, data_f0_out(159) => \data_f0_out[159]\, 
        data_f0_out(158) => \data_f0_out[158]\, data_f0_out(157)
         => \data_f0_out[157]\, data_f0_out(156) => 
        \data_f0_out[156]\, data_f0_out(155) => 
        \data_f0_out[155]\, data_f0_out(154) => 
        \data_f0_out[154]\, data_f0_out(153) => 
        \data_f0_out[153]\, data_f0_out(152) => 
        \data_f0_out[152]\, data_f0_out(151) => 
        \data_f0_out[151]\, data_f0_out(150) => 
        \data_f0_out[150]\, data_f0_out(149) => 
        \data_f0_out[149]\, data_f0_out(148) => 
        \data_f0_out[148]\, data_f0_out(147) => 
        \data_f0_out[147]\, data_f0_out(146) => 
        \data_f0_out[146]\, data_f0_out(145) => 
        \data_f0_out[145]\, data_f0_out(144) => 
        \data_f0_out[144]\, data_f0_out(143) => 
        \data_f0_out[143]\, data_f0_out(142) => 
        \data_f0_out[142]\, data_f0_out(141) => 
        \data_f0_out[141]\, data_f0_out(140) => 
        \data_f0_out[140]\, data_f0_out(139) => 
        \data_f0_out[139]\, data_f0_out(138) => 
        \data_f0_out[138]\, data_f0_out(137) => 
        \data_f0_out[137]\, data_f0_out(136) => 
        \data_f0_out[136]\, data_f0_out(135) => 
        \data_f0_out[135]\, data_f0_out(134) => 
        \data_f0_out[134]\, data_f0_out(133) => 
        \data_f0_out[133]\, data_f0_out(132) => 
        \data_f0_out[132]\, data_f0_out(131) => 
        \data_f0_out[131]\, data_f0_out(130) => 
        \data_f0_out[130]\, data_f0_out(129) => 
        \data_f0_out[129]\, data_f0_out(128) => 
        \data_f0_out[128]\, data_f0_out(127) => 
        \data_f0_out[127]\, data_f0_out(126) => 
        \data_f0_out[126]\, data_f0_out(125) => 
        \data_f0_out[125]\, data_f0_out(124) => 
        \data_f0_out[124]\, data_f0_out(123) => 
        \data_f0_out[123]\, data_f0_out(122) => 
        \data_f0_out[122]\, data_f0_out(121) => 
        \data_f0_out[121]\, data_f0_out(120) => 
        \data_f0_out[120]\, data_f0_out(119) => 
        \data_f0_out[119]\, data_f0_out(118) => 
        \data_f0_out[118]\, data_f0_out(117) => 
        \data_f0_out[117]\, data_f0_out(116) => 
        \data_f0_out[116]\, data_f0_out(115) => 
        \data_f0_out[115]\, data_f0_out(114) => 
        \data_f0_out[114]\, data_f0_out(113) => 
        \data_f0_out[113]\, data_f0_out(112) => 
        \data_f0_out[112]\, data_f0_out(111) => 
        \data_f0_out[111]\, data_f0_out(110) => 
        \data_f0_out[110]\, data_f0_out(109) => 
        \data_f0_out[109]\, data_f0_out(108) => 
        \data_f0_out[108]\, data_f0_out(107) => 
        \data_f0_out[107]\, data_f0_out(106) => 
        \data_f0_out[106]\, data_f0_out(105) => 
        \data_f0_out[105]\, data_f0_out(104) => 
        \data_f0_out[104]\, data_f0_out(103) => 
        \data_f0_out[103]\, data_f0_out(102) => 
        \data_f0_out[102]\, data_f0_out(101) => 
        \data_f0_out[101]\, data_f0_out(100) => 
        \data_f0_out[100]\, data_f0_out(99) => \data_f0_out[99]\, 
        data_f0_out(98) => \data_f0_out[98]\, data_f0_out(97) => 
        \data_f0_out[97]\, data_f0_out(96) => \data_f0_out[96]\, 
        data_f0_out(95) => \data_f0_out[95]\, data_f0_out(94) => 
        \data_f0_out[94]\, data_f0_out(93) => \data_f0_out[93]\, 
        data_f0_out(92) => \data_f0_out[92]\, data_f0_out(91) => 
        \data_f0_out[91]\, data_f0_out(90) => \data_f0_out[90]\, 
        data_f0_out(89) => \data_f0_out[89]\, data_f0_out(88) => 
        \data_f0_out[88]\, data_f0_out(87) => \data_f0_out[87]\, 
        data_f0_out(86) => \data_f0_out[86]\, data_f0_out(85) => 
        \data_f0_out[85]\, data_f0_out(84) => \data_f0_out[84]\, 
        data_f0_out(83) => \data_f0_out[83]\, data_f0_out(82) => 
        \data_f0_out[82]\, data_f0_out(81) => \data_f0_out[81]\, 
        data_f0_out(80) => \data_f0_out[80]\, data_f0_out(79) => 
        \data_f0_out[79]\, data_f0_out(78) => \data_f0_out[78]\, 
        data_f0_out(77) => \data_f0_out[77]\, data_f0_out(76) => 
        \data_f0_out[76]\, data_f0_out(75) => \data_f0_out[75]\, 
        data_f0_out(74) => \data_f0_out[74]\, data_f0_out(73) => 
        \data_f0_out[73]\, data_f0_out(72) => \data_f0_out[72]\, 
        data_f0_out(71) => \data_f0_out[71]\, data_f0_out(70) => 
        \data_f0_out[70]\, data_f0_out(69) => \data_f0_out[69]\, 
        data_f0_out(68) => \data_f0_out[68]\, data_f0_out(67) => 
        \data_f0_out[67]\, data_f0_out(66) => \data_f0_out[66]\, 
        data_f0_out(65) => \data_f0_out[65]\, data_f0_out(64) => 
        \data_f0_out[64]\, valid_out_i(1) => \valid_out_i[1]\, 
        ready_i_0(3) => \ready_i_0[3]\, ready_i_0(2) => 
        \ready_i_0[2]\, ready_i_0(1) => \ready_i_0[1]\, 
        ready_i_0(0) => \ready_i_0[0]\, valid_out_3 => 
        \valid_out[3]\, valid_out_2 => \valid_out[2]\, 
        valid_out_0 => \valid_out[0]\, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Downsampling_8_16_4 is

    port( sample_f0_0                   : out   std_logic;
          sample_f0_1                   : out   std_logic;
          sample_f0_2                   : out   std_logic;
          sample_f0_3                   : out   std_logic;
          sample_f0_4                   : out   std_logic;
          sample_f0_5                   : out   std_logic;
          sample_f0_6                   : out   std_logic;
          sample_f0_7                   : out   std_logic;
          sample_f0_8                   : out   std_logic;
          sample_f0_9                   : out   std_logic;
          sample_f0_10                  : out   std_logic;
          sample_f0_11                  : out   std_logic;
          sample_f0_12                  : out   std_logic;
          sample_f0_13                  : out   std_logic;
          sample_f0_14                  : out   std_logic;
          sample_f0_15                  : out   std_logic;
          sample_f0_32                  : out   std_logic;
          sample_f0_33                  : out   std_logic;
          sample_f0_34                  : out   std_logic;
          sample_f0_35                  : out   std_logic;
          sample_f0_36                  : out   std_logic;
          sample_f0_37                  : out   std_logic;
          sample_f0_38                  : out   std_logic;
          sample_f0_39                  : out   std_logic;
          sample_f0_40                  : out   std_logic;
          sample_f0_41                  : out   std_logic;
          sample_f0_42                  : out   std_logic;
          sample_f0_43                  : out   std_logic;
          sample_f0_44                  : out   std_logic;
          sample_f0_45                  : out   std_logic;
          sample_f0_46                  : out   std_logic;
          sample_f0_47                  : out   std_logic;
          sample_f0_48                  : out   std_logic;
          sample_f0_49                  : out   std_logic;
          sample_f0_50                  : out   std_logic;
          sample_f0_51                  : out   std_logic;
          sample_f0_52                  : out   std_logic;
          sample_f0_53                  : out   std_logic;
          sample_f0_54                  : out   std_logic;
          sample_f0_55                  : out   std_logic;
          sample_f0_56                  : out   std_logic;
          sample_f0_57                  : out   std_logic;
          sample_f0_58                  : out   std_logic;
          sample_f0_59                  : out   std_logic;
          sample_f0_60                  : out   std_logic;
          sample_f0_61                  : out   std_logic;
          sample_f0_62                  : out   std_logic;
          sample_f0_63                  : out   std_logic;
          sample_data_shaping_out_0     : in    std_logic;
          sample_data_shaping_out_1     : in    std_logic;
          sample_data_shaping_out_2     : in    std_logic;
          sample_data_shaping_out_3     : in    std_logic;
          sample_data_shaping_out_4     : in    std_logic;
          sample_data_shaping_out_5     : in    std_logic;
          sample_data_shaping_out_6     : in    std_logic;
          sample_data_shaping_out_7     : in    std_logic;
          sample_data_shaping_out_8     : in    std_logic;
          sample_data_shaping_out_9     : in    std_logic;
          sample_data_shaping_out_10    : in    std_logic;
          sample_data_shaping_out_11    : in    std_logic;
          sample_data_shaping_out_12    : in    std_logic;
          sample_data_shaping_out_13    : in    std_logic;
          sample_data_shaping_out_14    : in    std_logic;
          sample_data_shaping_out_15    : in    std_logic;
          sample_data_shaping_out_18    : in    std_logic;
          sample_data_shaping_out_19    : in    std_logic;
          sample_data_shaping_out_20    : in    std_logic;
          sample_data_shaping_out_21    : in    std_logic;
          sample_data_shaping_out_22    : in    std_logic;
          sample_data_shaping_out_23    : in    std_logic;
          sample_data_shaping_out_24    : in    std_logic;
          sample_data_shaping_out_25    : in    std_logic;
          sample_data_shaping_out_26    : in    std_logic;
          sample_data_shaping_out_27    : in    std_logic;
          sample_data_shaping_out_28    : in    std_logic;
          sample_data_shaping_out_29    : in    std_logic;
          sample_data_shaping_out_30    : in    std_logic;
          sample_data_shaping_out_31    : in    std_logic;
          sample_data_shaping_out_32    : in    std_logic;
          sample_data_shaping_out_33    : in    std_logic;
          sample_data_shaping_out_36    : in    std_logic;
          sample_data_shaping_out_37    : in    std_logic;
          sample_data_shaping_out_38    : in    std_logic;
          sample_data_shaping_out_39    : in    std_logic;
          sample_data_shaping_out_40    : in    std_logic;
          sample_data_shaping_out_41    : in    std_logic;
          sample_data_shaping_out_42    : in    std_logic;
          sample_data_shaping_out_43    : in    std_logic;
          sample_data_shaping_out_44    : in    std_logic;
          sample_data_shaping_out_45    : in    std_logic;
          sample_data_shaping_out_46    : in    std_logic;
          sample_data_shaping_out_47    : in    std_logic;
          sample_data_shaping_out_48    : in    std_logic;
          sample_data_shaping_out_49    : in    std_logic;
          sample_data_shaping_out_50    : in    std_logic;
          sample_data_shaping_out_51    : in    std_logic;
          sample_data_shaping_out_54    : in    std_logic;
          sample_data_shaping_out_55    : in    std_logic;
          sample_data_shaping_out_56    : in    std_logic;
          sample_data_shaping_out_57    : in    std_logic;
          sample_data_shaping_out_58    : in    std_logic;
          sample_data_shaping_out_59    : in    std_logic;
          sample_data_shaping_out_60    : in    std_logic;
          sample_data_shaping_out_61    : in    std_logic;
          sample_data_shaping_out_62    : in    std_logic;
          sample_data_shaping_out_63    : in    std_logic;
          sample_data_shaping_out_64    : in    std_logic;
          sample_data_shaping_out_65    : in    std_logic;
          sample_data_shaping_out_66    : in    std_logic;
          sample_data_shaping_out_67    : in    std_logic;
          sample_data_shaping_out_68    : in    std_logic;
          sample_data_shaping_out_69    : in    std_logic;
          sample_data_shaping_out_90    : in    std_logic;
          sample_data_shaping_out_91    : in    std_logic;
          sample_data_shaping_out_92    : in    std_logic;
          sample_data_shaping_out_93    : in    std_logic;
          sample_data_shaping_out_94    : in    std_logic;
          sample_data_shaping_out_95    : in    std_logic;
          sample_data_shaping_out_96    : in    std_logic;
          sample_data_shaping_out_97    : in    std_logic;
          sample_data_shaping_out_98    : in    std_logic;
          sample_data_shaping_out_99    : in    std_logic;
          sample_data_shaping_out_100   : in    std_logic;
          sample_data_shaping_out_101   : in    std_logic;
          sample_data_shaping_out_102   : in    std_logic;
          sample_data_shaping_out_103   : in    std_logic;
          sample_data_shaping_out_104   : in    std_logic;
          sample_data_shaping_out_105   : in    std_logic;
          sample_data_shaping_out_108   : in    std_logic;
          sample_data_shaping_out_109   : in    std_logic;
          sample_data_shaping_out_110   : in    std_logic;
          sample_data_shaping_out_111   : in    std_logic;
          sample_data_shaping_out_112   : in    std_logic;
          sample_data_shaping_out_113   : in    std_logic;
          sample_data_shaping_out_114   : in    std_logic;
          sample_data_shaping_out_115   : in    std_logic;
          sample_data_shaping_out_116   : in    std_logic;
          sample_data_shaping_out_117   : in    std_logic;
          sample_data_shaping_out_118   : in    std_logic;
          sample_data_shaping_out_119   : in    std_logic;
          sample_data_shaping_out_120   : in    std_logic;
          sample_data_shaping_out_121   : in    std_logic;
          sample_data_shaping_out_122   : in    std_logic;
          sample_data_shaping_out_123   : in    std_logic;
          sample_data_shaping_out_126   : in    std_logic;
          sample_data_shaping_out_127   : in    std_logic;
          sample_data_shaping_out_128   : in    std_logic;
          sample_data_shaping_out_129   : in    std_logic;
          sample_data_shaping_out_130   : in    std_logic;
          sample_data_shaping_out_131   : in    std_logic;
          sample_data_shaping_out_132   : in    std_logic;
          sample_data_shaping_out_133   : in    std_logic;
          sample_data_shaping_out_134   : in    std_logic;
          sample_data_shaping_out_135   : in    std_logic;
          sample_data_shaping_out_136   : in    std_logic;
          sample_data_shaping_out_137   : in    std_logic;
          sample_data_shaping_out_138   : in    std_logic;
          sample_data_shaping_out_139   : in    std_logic;
          sample_data_shaping_out_140   : in    std_logic;
          sample_data_shaping_out_141   : in    std_logic;
          sample_f0_wdata_95            : out   std_logic;
          sample_f0_wdata_94            : out   std_logic;
          sample_f0_wdata_93            : out   std_logic;
          sample_f0_wdata_92            : out   std_logic;
          sample_f0_wdata_91            : out   std_logic;
          sample_f0_wdata_90            : out   std_logic;
          sample_f0_wdata_89            : out   std_logic;
          sample_f0_wdata_88            : out   std_logic;
          sample_f0_wdata_87            : out   std_logic;
          sample_f0_wdata_86            : out   std_logic;
          sample_f0_wdata_85            : out   std_logic;
          sample_f0_wdata_84            : out   std_logic;
          sample_f0_wdata_83            : out   std_logic;
          sample_f0_wdata_82            : out   std_logic;
          sample_f0_wdata_81            : out   std_logic;
          sample_f0_wdata_80            : out   std_logic;
          sample_f0_wdata_79            : out   std_logic;
          sample_f0_wdata_78            : out   std_logic;
          sample_f0_wdata_77            : out   std_logic;
          sample_f0_wdata_76            : out   std_logic;
          sample_f0_wdata_75            : out   std_logic;
          sample_f0_wdata_74            : out   std_logic;
          sample_f0_wdata_73            : out   std_logic;
          sample_f0_wdata_72            : out   std_logic;
          sample_f0_wdata_71            : out   std_logic;
          sample_f0_wdata_70            : out   std_logic;
          sample_f0_wdata_69            : out   std_logic;
          sample_f0_wdata_68            : out   std_logic;
          sample_f0_wdata_67            : out   std_logic;
          sample_f0_wdata_66            : out   std_logic;
          sample_f0_wdata_65            : out   std_logic;
          sample_f0_wdata_64            : out   std_logic;
          sample_f0_wdata_63            : out   std_logic;
          sample_f0_wdata_62            : out   std_logic;
          sample_f0_wdata_61            : out   std_logic;
          sample_f0_wdata_60            : out   std_logic;
          sample_f0_wdata_59            : out   std_logic;
          sample_f0_wdata_58            : out   std_logic;
          sample_f0_wdata_57            : out   std_logic;
          sample_f0_wdata_56            : out   std_logic;
          sample_f0_wdata_55            : out   std_logic;
          sample_f0_wdata_54            : out   std_logic;
          sample_f0_wdata_53            : out   std_logic;
          sample_f0_wdata_52            : out   std_logic;
          sample_f0_wdata_51            : out   std_logic;
          sample_f0_wdata_50            : out   std_logic;
          sample_f0_wdata_49            : out   std_logic;
          sample_f0_wdata_48            : out   std_logic;
          sample_f0_wdata_15            : out   std_logic;
          sample_f0_wdata_14            : out   std_logic;
          sample_f0_wdata_13            : out   std_logic;
          sample_f0_wdata_12            : out   std_logic;
          sample_f0_wdata_11            : out   std_logic;
          sample_f0_wdata_10            : out   std_logic;
          sample_f0_wdata_9             : out   std_logic;
          sample_f0_wdata_8             : out   std_logic;
          sample_f0_wdata_7             : out   std_logic;
          sample_f0_wdata_6             : out   std_logic;
          sample_f0_wdata_5             : out   std_logic;
          sample_f0_wdata_4             : out   std_logic;
          sample_f0_wdata_3             : out   std_logic;
          sample_f0_wdata_2             : out   std_logic;
          sample_f0_wdata_1             : out   std_logic;
          sample_f0_wdata_0             : out   std_logic;
          sample_data_shaping_out_val   : in    std_logic;
          sample_f0_val                 : out   std_logic;
          sample_data_shaping_out_val_0 : in    std_logic;
          sample_f0_val_0               : out   std_logic;
          HRESETn_c                     : in    std_logic;
          HCLK_c                        : in    std_logic;
          sample_f0_val_1               : out   std_logic
        );

end Downsampling_8_16_4;

architecture DEF_ARCH of Downsampling_8_16_4 is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal sample_out_val_19, sample_out_0_sqmuxa_3, 
        un14_sample_in_val_0, sample_out_0_sqmuxa_2, 
        sample_out_0_sqmuxa_1, sample_out_0_sqmuxa_0, 
        un14_sample_in_val_23, un14_sample_in_val_22, 
        un14_sample_in_val_24, N_137, \counter[1]_net_1\, 
        \counter[0]_net_1\, N_129, \counter[3]_net_1\, 
        \DWACT_FDEC_E[0]\, N_106, \counter[8]_net_1\, 
        \DWACT_FDEC_E[4]\, N_91, \DWACT_FDEC_E[7]\, 
        \DWACT_FDEC_E[6]\, un14_sample_in_val_15, 
        un14_sample_in_val_14, un14_sample_in_val_20, 
        un14_sample_in_val_9, un14_sample_in_val_8, 
        un14_sample_in_val_19, un14_sample_in_val_5, 
        un14_sample_in_val_4, un14_sample_in_val_17, 
        un14_sample_in_val_13, \counter[24]_net_1\, 
        un14_sample_in_val_11, \counter[15]_net_1\, 
        \counter[12]_net_1\, un14_sample_in_val_7, 
        \counter[22]_net_1\, \counter[19]_net_1\, 
        un14_sample_in_val_3, \counter[23]_net_1\, 
        \counter[20]_net_1\, un14_sample_in_val_1, 
        \counter[11]_net_1\, \counter[27]_net_1\, 
        \counter[18]_net_1\, \counter[21]_net_1\, 
        \counter[9]_net_1\, \counter[4]_net_1\, 
        \counter[6]_net_1\, \counter[25]_net_1\, 
        \counter[2]_net_1\, \counter[13]_net_1\, 
        \counter[16]_net_1\, \counter[7]_net_1\, 
        \counter[10]_net_1\, \counter[26]_net_1\, 
        \counter[5]_net_1\, \counter[14]_net_1\, 
        \counter[17]_net_1\, un14_sample_in_val, 
        sample_out_0_sqmuxa, \counter_4[2]\, I_9, \counter_4[3]\, 
        I_13, \counter_4[4]\, I_20, \counter_4[5]\, I_24, 
        \counter_4[6]\, I_31_0, \counter_4[7]\, I_38, 
        \counter_4[8]\, I_45, \counter_4[9]\, I_52, 
        \counter_4[10]\, I_56, \counter_4[11]\, I_66, 
        \counter_4[12]\, I_73, \counter_4[13]\, I_77, 
        \counter_4[14]\, I_84, \counter_4[15]\, I_91, 
        \counter_4[16]\, I_98, \counter_4[17]\, I_105, 
        \counter_4[18]\, I_115, \counter_4[19]\, I_122, 
        \counter_4[20]\, I_129, \counter_4[21]\, I_136, 
        \counter_4[22]\, I_143, \counter_4[23]\, I_156, 
        \counter_4[24]\, I_166, \counter_4[25]\, I_173, 
        \counter_4[26]\, I_186, \counter_4[27]\, I_196, I_4, I_5, 
        N_4, \DWACT_FDEC_E[29]\, \DWACT_FDEC_E[30]\, 
        \DWACT_FDEC_E[23]\, \DWACT_FDEC_E[15]\, 
        \DWACT_FDEC_E[17]\, \DWACT_FDEC_E[22]\, N_11, 
        \DWACT_FDEC_E[21]\, \DWACT_FDEC_E[9]\, \DWACT_FDEC_E[12]\, 
        \DWACT_FDEC_E[20]\, N_20, \DWACT_FDEC_E[13]\, 
        \DWACT_FDEC_E[19]\, N_25, \DWACT_FDEC_E[18]\, N_32, 
        \DWACT_FDEC_E[33]\, \DWACT_FDEC_E[34]\, \DWACT_FDEC_E[2]\, 
        \DWACT_FDEC_E[5]\, N_41, \DWACT_FDEC_E[28]\, 
        \DWACT_FDEC_E[16]\, N_46, N_51, \DWACT_FDEC_E[14]\, N_56, 
        N_61, \DWACT_FDEC_E[10]\, N_68, \DWACT_FDEC_E[11]\, N_73, 
        N_78, N_83, \DWACT_FDEC_E[8]\, N_88, N_96, N_103, 
        \DWACT_FDEC_E[3]\, N_111, N_116, N_121, \DWACT_FDEC_E[1]\, 
        N_126, N_134, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \counter[19]\ : DFN1E1C0
      port map(D => \counter_4[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[19]_net_1\);
    
    \sample_out[125]\ : DFN1E1
      port map(D => sample_data_shaping_out_139, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_2);
    
    \sample_out[102]\ : DFN1E1
      port map(D => sample_data_shaping_out_114, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_54);
    
    \sample_out[122]\ : DFN1E1
      port map(D => sample_data_shaping_out_136, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_5);
    
    \sample_out[22]\ : DFN1E1
      port map(D => sample_data_shaping_out_24, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_73);
    
    \sample_out[101]\ : DFN1E1
      port map(D => sample_data_shaping_out_113, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_53);
    
    \sample_out[20]\ : DFN1E1
      port map(D => sample_data_shaping_out_22, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_75);
    
    \sample_out[13]\ : DFN1E1
      port map(D => sample_data_shaping_out_13, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_82);
    
    \sample_out[1]\ : DFN1E1
      port map(D => sample_data_shaping_out_1, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_94);
    
    \sample_out[19]\ : DFN1E1
      port map(D => sample_data_shaping_out_21, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_76);
    
    un3_counter_I_142 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[16]\, Y => N_41);
    
    \sample_out[61]\ : DFN1E1
      port map(D => sample_data_shaping_out_67, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_13);
    
    \sample_out[121]\ : DFN1E1
      port map(D => sample_data_shaping_out_135, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_6);
    
    \sample_out[38]\ : DFN1E1
      port map(D => sample_data_shaping_out_42, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_57);
    
    un3_counter_I_27 : OR2
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        Y => \DWACT_FDEC_E[1]\);
    
    \sample_out[95]\ : DFN1E1
      port map(D => sample_data_shaping_out_105, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_47);
    
    \counter_RNO[11]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_66, Y => 
        \counter_4[11]\);
    
    \counter_RNIHDLE1[10]\ : NOR3B
      port map(A => sample_data_shaping_out_val_0, B => HRESETn_c, 
        C => un14_sample_in_val_0, Y => sample_out_0_sqmuxa_1);
    
    \sample_out[104]\ : DFN1E1
      port map(D => sample_data_shaping_out_116, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_56);
    
    \sample_out[34]\ : DFN1E1
      port map(D => sample_data_shaping_out_38, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_61);
    
    un3_counter_I_4 : INV
      port map(A => \counter[0]_net_1\, Y => I_4);
    
    \sample_out[124]\ : DFN1E1
      port map(D => sample_data_shaping_out_138, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_3);
    
    \counter[11]\ : DFN1E1C0
      port map(D => \counter_4[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[11]_net_1\);
    
    un3_counter_I_94 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, Y
         => \DWACT_FDEC_E[10]\);
    
    \counter_RNI0L371[10]\ : OR3C
      port map(A => un14_sample_in_val_23, B => 
        un14_sample_in_val_22, C => un14_sample_in_val_24, Y => 
        un14_sample_in_val_0);
    
    \sample_out[97]\ : DFN1E1
      port map(D => sample_data_shaping_out_109, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_49);
    
    un3_counter_I_186 : XNOR2
      port map(A => N_11, B => \counter[26]_net_1\, Y => I_186);
    
    \sample_out[108]\ : DFN1E1
      port map(D => sample_data_shaping_out_120, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_60);
    
    \counter_RNO[15]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_91, Y => 
        \counter_4[15]\);
    
    un3_counter_I_108 : OR3
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        C => \counter[17]_net_1\, Y => \DWACT_FDEC_E[12]\);
    
    un3_counter_I_121 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \counter[18]_net_1\, Y => N_56);
    
    \sample_out[51]\ : DFN1E1
      port map(D => sample_data_shaping_out_57, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_3);
    
    \sample_out[56]\ : DFN1E1
      port map(D => sample_data_shaping_out_62, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_8);
    
    un3_counter_I_176 : OR2
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        Y => \DWACT_FDEC_E[20]\);
    
    \sample_out[0]\ : DFN1E1
      port map(D => sample_data_shaping_out_0, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_95);
    
    \counter_RNO[7]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_38, Y => 
        \counter_4[7]\);
    
    \counter[6]\ : DFN1E1C0
      port map(D => \counter_4[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[6]_net_1\);
    
    un3_counter_I_48 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => \DWACT_FDEC_E[4]\);
    
    un3_counter_I_114 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[10]\, 
        C => \DWACT_FDEC_E[12]\, Y => N_61);
    
    \counter[21]\ : DFN1E1C0
      port map(D => \counter_4[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[21]_net_1\);
    
    un3_counter_I_13 : XNOR2
      port map(A => N_134, B => \counter[3]_net_1\, Y => I_13);
    
    \sample_out[81]\ : DFN1E1
      port map(D => sample_data_shaping_out_91, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_33);
    
    \sample_out[86]\ : DFN1E1
      port map(D => sample_data_shaping_out_96, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_38);
    
    \counter[3]\ : DFN1E1C0
      port map(D => \counter_4[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[3]_net_1\);
    
    \counter[2]\ : DFN1E1C0
      port map(D => \counter_4[2]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[2]_net_1\);
    
    un3_counter_I_73 : XNOR2
      port map(A => N_91, B => \counter[12]_net_1\, Y => I_73);
    
    \counter_RNO[8]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_45, Y => 
        \counter_4[8]\);
    
    \counter_RNO[13]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_77, Y => 
        \counter_4[13]\);
    
    un3_counter_I_52 : XNOR2
      port map(A => N_106, B => \counter[9]_net_1\, Y => I_52);
    
    \counter_RNIKF54[20]\ : NOR3A
      port map(A => un14_sample_in_val_3, B => 
        \counter[23]_net_1\, C => \counter[20]_net_1\, Y => 
        un14_sample_in_val_15);
    
    \sample_out[12]\ : DFN1E1
      port map(D => sample_data_shaping_out_12, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_83);
    
    \sample_out[10]\ : DFN1E1
      port map(D => sample_data_shaping_out_10, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_85);
    
    \sample_out[45]\ : DFN1E1
      port map(D => sample_data_shaping_out_49, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_50);
    
    \counter_RNO[12]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_73, Y => 
        \counter_4[12]\);
    
    \sample_out[33]\ : DFN1E1
      port map(D => sample_data_shaping_out_37, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_62);
    
    \sample_out[39]\ : DFN1E1
      port map(D => sample_data_shaping_out_43, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_56);
    
    \counter[17]\ : DFN1E1C0
      port map(D => \counter_4[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[17]_net_1\);
    
    un3_counter_I_41 : OR2
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        Y => \DWACT_FDEC_E[3]\);
    
    un3_counter_I_159 : OR3
      port map(A => \counter[21]_net_1\, B => \counter[22]_net_1\, 
        C => \counter[23]_net_1\, Y => \DWACT_FDEC_E[17]\);
    
    \counter[4]\ : DFN1E1C0
      port map(D => \counter_4[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[4]_net_1\);
    
    un3_counter_I_5 : XNOR2
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        Y => I_5);
    
    un3_counter_I_125 : OR2
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        Y => \DWACT_FDEC_E[14]\);
    
    \counter[10]\ : DFN1E1C0
      port map(D => \counter_4[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[10]_net_1\);
    
    \sample_out[5]\ : DFN1E1
      port map(D => sample_data_shaping_out_5, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_wdata_90);
    
    \sample_out[47]\ : DFN1E1
      port map(D => sample_data_shaping_out_51, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_wdata_48);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter[13]\ : DFN1E1C0
      port map(D => \counter_4[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[13]_net_1\);
    
    un3_counter_I_62 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[6]\);
    
    \counter_RNILSE[14]\ : NOR2
      port map(A => \counter[14]_net_1\, B => \counter[17]_net_1\, 
        Y => un14_sample_in_val_1);
    
    un3_counter_I_139 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        Y => \DWACT_FDEC_E[16]\);
    
    \sample_out[115]\ : DFN1E1
      port map(D => sample_data_shaping_out_129, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_12);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sample_out[21]\ : DFN1E1
      port map(D => sample_data_shaping_out_23, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_74);
    
    \counter[12]\ : DFN1E1C0
      port map(D => \counter_4[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[12]_net_1\);
    
    \sample_out[26]\ : DFN1E1
      port map(D => sample_data_shaping_out_28, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_69);
    
    \counter_RNIB507[3]\ : NOR2
      port map(A => \counter[3]_net_1\, B => \counter[0]_net_1\, 
        Y => un14_sample_in_val_13);
    
    \sample_out[2]\ : DFN1E1
      port map(D => sample_data_shaping_out_2, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_93);
    
    \sample_out[98]\ : DFN1E1
      port map(D => sample_data_shaping_out_110, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_50);
    
    \sample_out[112]\ : DFN1E1
      port map(D => sample_data_shaping_out_126, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_15);
    
    \counter_RNIHDLE1_1[10]\ : NOR3B
      port map(A => sample_data_shaping_out_val_0, B => HRESETn_c, 
        C => un14_sample_in_val_0, Y => sample_out_0_sqmuxa_0);
    
    \counter[27]\ : DFN1E1C0
      port map(D => \counter_4[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[27]_net_1\);
    
    un3_counter_I_111 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[28]\);
    
    \counter[20]\ : DFN1E1C0
      port map(D => \counter_4[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[20]_net_1\);
    
    \sample_out[94]\ : DFN1E1
      port map(D => sample_data_shaping_out_104, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_46);
    
    \sample_out[111]\ : DFN1E1
      port map(D => sample_data_shaping_out_123, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_63);
    
    un3_counter_I_166 : XNOR2
      port map(A => N_25, B => \counter[24]_net_1\, Y => I_166);
    
    \counter_RNO[17]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_105, Y => 
        \counter_4[17]\);
    
    \counter_RNII3CB1[10]\ : NOR2A
      port map(A => sample_data_shaping_out_val_0, B => 
        un14_sample_in_val_0, Y => sample_out_val_19);
    
    \counter[23]\ : DFN1E1C0
      port map(D => \counter_4[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[23]_net_1\);
    
    \counter_RNIGCTE[12]\ : NOR3C
      port map(A => un14_sample_in_val_9, B => 
        un14_sample_in_val_8, C => un14_sample_in_val_19, Y => 
        un14_sample_in_val_23);
    
    \counter_RNI8DT[27]\ : NOR3A
      port map(A => un14_sample_in_val_1, B => 
        \counter[11]_net_1\, C => \counter[27]_net_1\, Y => 
        un14_sample_in_val_14);
    
    un3_counter_I_149 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[34]\);
    
    \sample_out[55]\ : DFN1E1
      port map(D => sample_data_shaping_out_61, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_7);
    
    \counter[22]\ : DFN1E1C0
      port map(D => \counter_4[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[22]_net_1\);
    
    \counter[15]\ : DFN1E1C0
      port map(D => \counter_4[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[15]_net_1\);
    
    un3_counter_I_8 : OR2
      port map(A => \counter[1]_net_1\, B => \counter[0]_net_1\, 
        Y => N_137);
    
    un3_counter_I_185 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[21]\, Y => N_11);
    
    \sample_out[114]\ : DFN1E1
      port map(D => sample_data_shaping_out_128, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_13);
    
    un3_counter_I_196 : XNOR2
      port map(A => N_4, B => \counter[27]_net_1\, Y => I_196);
    
    \counter_RNIHDLE1_0[10]\ : NOR3B
      port map(A => sample_data_shaping_out_val_0, B => HRESETn_c, 
        C => un14_sample_in_val_0, Y => sample_out_0_sqmuxa_2);
    
    \sample_out[32]\ : DFN1E1
      port map(D => sample_data_shaping_out_36, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_63);
    
    un3_counter_I_51 : OR2
      port map(A => \counter[8]_net_1\, B => \DWACT_FDEC_E[4]\, Y
         => N_106);
    
    un3_counter_I_122 : XNOR2
      port map(A => N_56, B => \counter[19]_net_1\, Y => I_122);
    
    \sample_out[118]\ : DFN1E1
      port map(D => sample_data_shaping_out_132, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_9);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sample_out[57]\ : DFN1E1
      port map(D => sample_data_shaping_out_63, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_9);
    
    \sample_out[30]\ : DFN1E1
      port map(D => sample_data_shaping_out_32, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_65);
    
    \counter_RNO[14]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_84, Y => 
        \counter_4[14]\);
    
    \sample_out[85]\ : DFN1E1
      port map(D => sample_data_shaping_out_95, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_37);
    
    \counter_RNI51T[12]\ : NOR3A
      port map(A => un14_sample_in_val_11, B => 
        \counter[15]_net_1\, C => \counter[12]_net_1\, Y => 
        un14_sample_in_val_19);
    
    \counter[1]\ : DFN1E1C0
      port map(D => I_5, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_data_shaping_out_val, Q => \counter[1]_net_1\);
    
    \counter_RNO[26]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_186, Y => 
        \counter_4[26]\);
    
    \sample_out[4]\ : DFN1E1
      port map(D => sample_data_shaping_out_4, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_wdata_91);
    
    \counter_RNO[5]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_24, Y => 
        \counter_4[5]\);
    
    \sample_out[103]\ : DFN1E1
      port map(D => sample_data_shaping_out_115, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_55);
    
    \sample_out[100]\ : DFN1E1
      port map(D => sample_data_shaping_out_112, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_52);
    
    \counter[25]\ : DFN1E1C0
      port map(D => \counter_4[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[25]_net_1\);
    
    \sample_out[123]\ : DFN1E1
      port map(D => sample_data_shaping_out_137, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_4);
    
    \sample_out[120]\ : DFN1E1
      port map(D => sample_data_shaping_out_134, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_7);
    
    \counter_RNI0RM3[10]\ : NOR2
      port map(A => \counter[7]_net_1\, B => \counter[10]_net_1\, 
        Y => un14_sample_in_val_4);
    
    sample_out_val : DFN1C0
      port map(D => sample_out_val_19, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f0_val);
    
    \counter_RNO[3]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_13, Y => 
        \counter_4[3]\);
    
    \sample_out[87]\ : DFN1E1
      port map(D => sample_data_shaping_out_97, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_39);
    
    un3_counter_I_115 : XNOR2
      port map(A => N_61, B => \counter[18]_net_1\, Y => I_115);
    
    un3_counter_I_87 : OR3
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        C => \counter[14]_net_1\, Y => \DWACT_FDEC_E[9]\);
    
    un3_counter_I_173 : XNOR2
      port map(A => N_20, B => \counter[25]_net_1\, Y => I_173);
    
    \sample_out[48]\ : DFN1E1
      port map(D => sample_data_shaping_out_54, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_0);
    
    un3_counter_I_38 : XNOR2
      port map(A => N_116, B => \counter[7]_net_1\, Y => I_38);
    
    \sample_out[93]\ : DFN1E1
      port map(D => sample_data_shaping_out_103, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_45);
    
    \sample_out[11]\ : DFN1E1
      port map(D => sample_data_shaping_out_11, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_84);
    
    \sample_out[99]\ : DFN1E1
      port map(D => sample_data_shaping_out_111, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_51);
    
    \sample_out[16]\ : DFN1E1
      port map(D => sample_data_shaping_out_18, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_79);
    
    \counter[5]\ : DFN1E1C0
      port map(D => \counter_4[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[5]_net_1\);
    
    \counter_RNIAGNA[24]\ : NOR3A
      port map(A => un14_sample_in_val_13, B => 
        \counter[1]_net_1\, C => \counter[24]_net_1\, Y => 
        un14_sample_in_val_20);
    
    \sample_out[44]\ : DFN1E1
      port map(D => sample_data_shaping_out_48, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_51);
    
    \counter_RNIP507[8]\ : NOR2
      port map(A => \counter[8]_net_1\, B => \counter[9]_net_1\, 
        Y => un14_sample_in_val_9);
    
    \counter_RNIJKE[13]\ : NOR2
      port map(A => \counter[13]_net_1\, B => \counter[16]_net_1\, 
        Y => un14_sample_in_val_5);
    
    un3_counter_I_37 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \counter[6]_net_1\, Y => N_116);
    
    \counter_RNINB64[22]\ : NOR3A
      port map(A => un14_sample_in_val_7, B => 
        \counter[22]_net_1\, C => \counter[19]_net_1\, Y => 
        un14_sample_in_val_17);
    
    \counter_RNO[10]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_56, Y => 
        \counter_4[10]\);
    
    un3_counter_I_9 : XNOR2
      port map(A => N_137, B => \counter[2]_net_1\, Y => I_9);
    
    \counter_RNO[21]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_136, Y => 
        \counter_4[21]\);
    
    un3_counter_I_20 : XNOR2
      port map(A => N_129, B => \counter[4]_net_1\, Y => I_20);
    
    un3_counter_I_182 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[30]\);
    
    \sample_out[25]\ : DFN1E1
      port map(D => sample_data_shaping_out_27, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_70);
    
    un3_counter_I_56 : XNOR2
      port map(A => N_103, B => \counter[10]_net_1\, Y => I_56);
    
    \counter[16]\ : DFN1E1C0
      port map(D => \counter_4[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[16]_net_1\);
    
    \counter_RNO[25]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_173, Y => 
        \counter_4[25]\);
    
    un3_counter_I_172 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[19]\, Y => N_20);
    
    un3_counter_I_104 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \DWACT_FDEC_E[11]\, Y => N_68);
    
    un3_counter_I_31 : XNOR2
      port map(A => N_121, B => \counter[6]_net_1\, Y => I_31_0);
    
    un3_counter_I_98 : XNOR2
      port map(A => N_73, B => \counter[16]_net_1\, Y => I_98);
    
    \counter_RNIHDLE1_3[10]\ : NOR3B
      port map(A => sample_data_shaping_out_val_0, B => HRESETn_c, 
        C => un14_sample_in_val_0, Y => sample_out_0_sqmuxa);
    
    un3_counter_I_23 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \counter[3]_net_1\, C
         => \counter[4]_net_1\, Y => N_126);
    
    \sample_out[27]\ : DFN1E1
      port map(D => sample_data_shaping_out_29, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_68);
    
    un3_counter_I_59 : OR3
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        C => \counter[8]_net_1\, Y => \DWACT_FDEC_E[5]\);
    
    un3_counter_I_12 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => N_134);
    
    \counter_RNO[6]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_31_0, Y => 
        \counter_4[6]\);
    
    un3_counter_I_165 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[18]\, Y => N_25);
    
    \counter_RNI6DQF[20]\ : NOR3C
      port map(A => un14_sample_in_val_15, B => 
        un14_sample_in_val_14, C => un14_sample_in_val_20, Y => 
        un14_sample_in_val_24);
    
    un3_counter_I_156 : XNOR2
      port map(A => N_32, B => \counter[23]_net_1\, Y => I_156);
    
    un3_counter_I_97 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \counter[15]_net_1\, Y => N_73);
    
    un3_counter_I_128 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[14]\, Y => N_51);
    
    un3_counter_I_72 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[6]\, Y
         => N_91);
    
    \sample_out[58]\ : DFN1E1
      port map(D => sample_data_shaping_out_64, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_10);
    
    \counter[26]\ : DFN1E1C0
      port map(D => \counter_4[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[26]_net_1\);
    
    un3_counter_I_66 : XNOR2
      port map(A => N_96, B => \counter[11]_net_1\, Y => I_66);
    
    \counter_RNO[23]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_156, Y => 
        \counter_4[23]\);
    
    \sample_out[54]\ : DFN1E1
      port map(D => sample_data_shaping_out_60, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_6);
    
    \sample_out[43]\ : DFN1E1
      port map(D => sample_data_shaping_out_47, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_52);
    
    \sample_out[49]\ : DFN1E1
      port map(D => sample_data_shaping_out_55, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_1);
    
    sample_out_val_0 : DFN1C0
      port map(D => sample_out_val_19, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f0_val_0);
    
    un3_counter_I_45 : XNOR2
      port map(A => N_111, B => \counter[8]_net_1\, Y => I_45);
    
    un3_counter_I_24 : XNOR2
      port map(A => N_126, B => \counter[5]_net_1\, Y => I_24);
    
    un3_counter_I_195 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[23]\, Y => N_4);
    
    \sample_out[92]\ : DFN1E1
      port map(D => sample_data_shaping_out_102, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_44);
    
    \counter[14]\ : DFN1E1C0
      port map(D => \counter_4[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[14]_net_1\);
    
    un3_counter_I_136 : XNOR2
      port map(A => N_46, B => \counter[21]_net_1\, Y => I_136);
    
    \sample_out[88]\ : DFN1E1
      port map(D => sample_data_shaping_out_98, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_40);
    
    \sample_out[90]\ : DFN1E1
      port map(D => sample_data_shaping_out_100, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_42);
    
    un3_counter_I_91 : XNOR2
      port map(A => N_78, B => \counter[15]_net_1\, Y => I_91);
    
    \counter_RNO[22]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_143, Y => 
        \counter_4[22]\);
    
    \sample_out[31]\ : DFN1E1
      port map(D => sample_data_shaping_out_33, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_64);
    
    \sample_out[36]\ : DFN1E1
      port map(D => sample_data_shaping_out_40, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_59);
    
    un3_counter_I_69 : OR3
      port map(A => \counter[9]_net_1\, B => \counter[10]_net_1\, 
        C => \counter[11]_net_1\, Y => \DWACT_FDEC_E[7]\);
    
    \sample_out[84]\ : DFN1E1
      port map(D => sample_data_shaping_out_94, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_36);
    
    \sample_out[63]\ : DFN1E1
      port map(D => sample_data_shaping_out_69, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_15);
    
    \counter_RNI5JN3[26]\ : NOR2
      port map(A => \counter[26]_net_1\, B => \counter[5]_net_1\, 
        Y => un14_sample_in_val_3);
    
    \sample_out[15]\ : DFN1E1
      port map(D => sample_data_shaping_out_15, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_80);
    
    un3_counter_I_129 : XNOR2
      port map(A => N_51, B => \counter[20]_net_1\, Y => I_129);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un3_counter_I_146 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        C => \counter[22]_net_1\, Y => \DWACT_FDEC_E[33]\);
    
    \counter[24]\ : DFN1E1C0
      port map(D => \counter_4[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[24]_net_1\);
    
    un3_counter_I_101 : OR2
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        Y => \DWACT_FDEC_E[11]\);
    
    \sample_out[113]\ : DFN1E1
      port map(D => sample_data_shaping_out_127, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_14);
    
    \sample_out[110]\ : DFN1E1
      port map(D => sample_data_shaping_out_122, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_62);
    
    \counter_RNO[4]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_20, Y => 
        \counter_4[4]\);
    
    un3_counter_I_162 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        Y => \DWACT_FDEC_E[18]\);
    
    \sample_out[106]\ : DFN1E1
      port map(D => sample_data_shaping_out_118, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_58);
    
    un3_counter_I_77 : XNOR2
      port map(A => N_88, B => \counter[13]_net_1\, Y => I_77);
    
    \sample_out[17]\ : DFN1E1
      port map(D => sample_data_shaping_out_19, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_78);
    
    \sample_out[107]\ : DFN1E1
      port map(D => sample_data_shaping_out_119, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_59);
    
    \counter_RNO[18]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_115, Y => 
        \counter_4[18]\);
    
    un3_counter_I_44 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => N_111);
    
    \sample_out[126]\ : DFN1E1
      port map(D => sample_data_shaping_out_140, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_1);
    
    \sample_out[127]\ : DFN1E1
      port map(D => sample_data_shaping_out_141, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_0);
    
    \counter_RNIKKE[21]\ : NOR2
      port map(A => \counter[18]_net_1\, B => \counter[21]_net_1\, 
        Y => un14_sample_in_val_11);
    
    \sample_out[53]\ : DFN1E1
      port map(D => sample_data_shaping_out_59, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_5);
    
    \sample_out[28]\ : DFN1E1
      port map(D => sample_data_shaping_out_30, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_67);
    
    \counter_RNO[27]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_196, Y => 
        \counter_4[27]\);
    
    \sample_out[59]\ : DFN1E1
      port map(D => sample_data_shaping_out_65, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_11);
    
    \sample_out[109]\ : DFN1E1
      port map(D => sample_data_shaping_out_121, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_61);
    
    un3_counter_I_192 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[22]\, Y => \DWACT_FDEC_E[23]\);
    
    \sample_out[24]\ : DFN1E1
      port map(D => sample_data_shaping_out_26, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_71);
    
    un3_counter_I_55 : OR3
      port map(A => \DWACT_FDEC_E[4]\, B => \counter[8]_net_1\, C
         => \counter[9]_net_1\, Y => N_103);
    
    \sample_out[42]\ : DFN1E1
      port map(D => sample_data_shaping_out_46, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_53);
    
    un3_counter_I_118 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[13]\);
    
    \sample_out[40]\ : DFN1E1
      port map(D => sample_data_shaping_out_44, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_55);
    
    \sample_out[83]\ : DFN1E1
      port map(D => sample_data_shaping_out_93, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_35);
    
    \sample_out[89]\ : DFN1E1
      port map(D => sample_data_shaping_out_99, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_41);
    
    un3_counter_I_189 : OR3
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        C => \counter[26]_net_1\, Y => \DWACT_FDEC_E[22]\);
    
    \counter_RNO[24]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_166, Y => 
        \counter_4[24]\);
    
    \counter[7]\ : DFN1E1C0
      port map(D => \counter_4[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[7]_net_1\);
    
    un3_counter_I_105 : XNOR2
      port map(A => N_68, B => \counter[17]_net_1\, Y => I_105);
    
    \sample_out[6]\ : DFN1E1
      port map(D => sample_data_shaping_out_6, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_wdata_89);
    
    un3_counter_I_155 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[33]\, Y => N_32);
    
    un3_counter_I_179 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[20]\, Y => \DWACT_FDEC_E[21]\);
    
    \sample_out[62]\ : DFN1E1
      port map(D => sample_data_shaping_out_68, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_14);
    
    \sample_out[60]\ : DFN1E1
      port map(D => sample_data_shaping_out_66, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_12);
    
    un3_counter_I_65 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \counter[9]_net_1\, C
         => \counter[10]_net_1\, Y => N_96);
    
    \sample_out[35]\ : DFN1E1
      port map(D => sample_data_shaping_out_39, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_60);
    
    \sample_out[91]\ : DFN1E1
      port map(D => sample_data_shaping_out_101, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_43);
    
    un3_counter_I_135 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[15]\, Y => N_46);
    
    \sample_out[96]\ : DFN1E1
      port map(D => sample_data_shaping_out_108, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_48);
    
    un3_counter_I_80 : OR2
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        Y => \DWACT_FDEC_E[8]\);
    
    \counter_RNII507[4]\ : NOR2
      port map(A => \counter[4]_net_1\, B => \counter[6]_net_1\, 
        Y => un14_sample_in_val_8);
    
    un3_counter_I_16 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[0]\);
    
    \counter_RNI1FN3[25]\ : NOR2
      port map(A => \counter[25]_net_1\, B => \counter[2]_net_1\, 
        Y => un14_sample_in_val_7);
    
    sample_out_val_1 : DFN1C0
      port map(D => sample_out_val_19, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f0_val_1);
    
    \counter_RNO[20]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_129, Y => 
        \counter_4[20]\);
    
    \sample_out[37]\ : DFN1E1
      port map(D => sample_data_shaping_out_41, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_58);
    
    \sample_out[23]\ : DFN1E1
      port map(D => sample_data_shaping_out_25, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_72);
    
    \sample_out[52]\ : DFN1E1
      port map(D => sample_data_shaping_out_58, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_4);
    
    \sample_out[29]\ : DFN1E1
      port map(D => sample_data_shaping_out_31, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_66);
    
    un3_counter_I_76 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \counter[12]_net_1\, Y => N_88);
    
    un3_counter_I_30 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[1]\, C
         => \counter[5]_net_1\, Y => N_121);
    
    \sample_out[50]\ : DFN1E1
      port map(D => sample_data_shaping_out_56, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_2);
    
    \sample_out[18]\ : DFN1E1
      port map(D => sample_data_shaping_out_20, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_77);
    
    \sample_out[9]\ : DFN1E1
      port map(D => sample_data_shaping_out_9, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_wdata_86);
    
    \sample_out[7]\ : DFN1E1
      port map(D => sample_data_shaping_out_7, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_wdata_88);
    
    un3_counter_I_83 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[8]\, Y => N_83);
    
    un3_counter_I_19 : OR2
      port map(A => \counter[3]_net_1\, B => \DWACT_FDEC_E[0]\, Y
         => N_129);
    
    \sample_out[14]\ : DFN1E1
      port map(D => sample_data_shaping_out_14, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_1, Q => sample_f0_wdata_81);
    
    \counter_RNIHDLE1_2[10]\ : NOR3B
      port map(A => sample_data_shaping_out_val_0, B => HRESETn_c, 
        C => un14_sample_in_val_0, Y => sample_out_0_sqmuxa_3);
    
    \sample_out[82]\ : DFN1E1
      port map(D => sample_data_shaping_out_92, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_34);
    
    \counter_RNO[2]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_9, Y => 
        \counter_4[2]\);
    
    \counter[9]\ : DFN1E1C0
      port map(D => \counter_4[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[9]_net_1\);
    
    \sample_out[80]\ : DFN1E1
      port map(D => sample_data_shaping_out_90, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_3, Q => sample_f0_32);
    
    \counter_RNO[19]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_122, Y => 
        \counter_4[19]\);
    
    \counter_RNIARB8[10]\ : NOR3C
      port map(A => un14_sample_in_val_5, B => 
        un14_sample_in_val_4, C => un14_sample_in_val_17, Y => 
        un14_sample_in_val_22);
    
    un3_counter_I_152 : OR3
      port map(A => \DWACT_FDEC_E[34]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[29]\);
    
    \counter_RNO[9]\ : NOR2B
      port map(A => un14_sample_in_val_0, B => I_52, Y => 
        \counter_4[9]\);
    
    \counter_RNI0L371_0[10]\ : OR3C
      port map(A => un14_sample_in_val_23, B => 
        un14_sample_in_val_22, C => un14_sample_in_val_24, Y => 
        un14_sample_in_val);
    
    \counter[8]\ : DFN1E1C0
      port map(D => \counter_4[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val, Q => 
        \counter[8]_net_1\);
    
    un3_counter_I_84 : XNOR2
      port map(A => N_83, B => \counter[14]_net_1\, Y => I_84);
    
    un3_counter_I_143 : XNOR2
      port map(A => N_41, B => \counter[22]_net_1\, Y => I_143);
    
    \sample_out[116]\ : DFN1E1
      port map(D => sample_data_shaping_out_130, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_11);
    
    \counter[18]\ : DFN1E1C0
      port map(D => \counter_4[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_data_shaping_out_val_0, Q => 
        \counter[18]_net_1\);
    
    \sample_out[117]\ : DFN1E1
      port map(D => sample_data_shaping_out_131, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_10);
    
    un3_counter_I_90 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[9]\, Y => N_78);
    
    un3_counter_I_169 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \counter[24]_net_1\, Y => \DWACT_FDEC_E[19]\);
    
    un3_counter_I_132 : OR3
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        C => \counter[20]_net_1\, Y => \DWACT_FDEC_E[15]\);
    
    \sample_out[8]\ : DFN1E1
      port map(D => sample_data_shaping_out_8, CLK => HCLK_c, E
         => sample_out_0_sqmuxa, Q => sample_f0_wdata_87);
    
    \sample_out[41]\ : DFN1E1
      port map(D => sample_data_shaping_out_45, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_54);
    
    \counter_RNO[16]\ : NOR2B
      port map(A => un14_sample_in_val, B => I_98, Y => 
        \counter_4[16]\);
    
    \counter[0]\ : DFN1E1C0
      port map(D => I_4, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_data_shaping_out_val_0, Q => \counter[0]_net_1\);
    
    \sample_out[46]\ : DFN1E1
      port map(D => sample_data_shaping_out_50, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_49);
    
    \sample_out[3]\ : DFN1E1
      port map(D => sample_data_shaping_out_3, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_2, Q => sample_f0_wdata_92);
    
    un3_counter_I_34 : OR3
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        C => \counter[5]_net_1\, Y => \DWACT_FDEC_E[2]\);
    
    \sample_out[105]\ : DFN1E1
      port map(D => sample_data_shaping_out_117, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_57);
    
    \sample_out[119]\ : DFN1E1
      port map(D => sample_data_shaping_out_133, CLK => HCLK_c, E
         => sample_out_0_sqmuxa_0, Q => sample_f0_wdata_8);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity Downsampling_8_16_6 is

    port( sample_f0_0           : in    std_logic;
          sample_f0_1           : in    std_logic;
          sample_f0_2           : in    std_logic;
          sample_f0_3           : in    std_logic;
          sample_f0_4           : in    std_logic;
          sample_f0_5           : in    std_logic;
          sample_f0_6           : in    std_logic;
          sample_f0_7           : in    std_logic;
          sample_f0_8           : in    std_logic;
          sample_f0_9           : in    std_logic;
          sample_f0_10          : in    std_logic;
          sample_f0_11          : in    std_logic;
          sample_f0_12          : in    std_logic;
          sample_f0_13          : in    std_logic;
          sample_f0_14          : in    std_logic;
          sample_f0_15          : in    std_logic;
          sample_f0_32          : in    std_logic;
          sample_f0_33          : in    std_logic;
          sample_f0_34          : in    std_logic;
          sample_f0_35          : in    std_logic;
          sample_f0_36          : in    std_logic;
          sample_f0_37          : in    std_logic;
          sample_f0_38          : in    std_logic;
          sample_f0_39          : in    std_logic;
          sample_f0_40          : in    std_logic;
          sample_f0_41          : in    std_logic;
          sample_f0_42          : in    std_logic;
          sample_f0_43          : in    std_logic;
          sample_f0_44          : in    std_logic;
          sample_f0_45          : in    std_logic;
          sample_f0_46          : in    std_logic;
          sample_f0_47          : in    std_logic;
          sample_f0_48          : in    std_logic;
          sample_f0_49          : in    std_logic;
          sample_f0_50          : in    std_logic;
          sample_f0_51          : in    std_logic;
          sample_f0_52          : in    std_logic;
          sample_f0_53          : in    std_logic;
          sample_f0_54          : in    std_logic;
          sample_f0_55          : in    std_logic;
          sample_f0_56          : in    std_logic;
          sample_f0_57          : in    std_logic;
          sample_f0_58          : in    std_logic;
          sample_f0_59          : in    std_logic;
          sample_f0_60          : in    std_logic;
          sample_f0_61          : in    std_logic;
          sample_f0_62          : in    std_logic;
          sample_f0_63          : in    std_logic;
          sample_f1_0           : out   std_logic;
          sample_f1_1           : out   std_logic;
          sample_f1_2           : out   std_logic;
          sample_f1_3           : out   std_logic;
          sample_f1_4           : out   std_logic;
          sample_f1_5           : out   std_logic;
          sample_f1_6           : out   std_logic;
          sample_f1_7           : out   std_logic;
          sample_f1_8           : out   std_logic;
          sample_f1_9           : out   std_logic;
          sample_f1_10          : out   std_logic;
          sample_f1_11          : out   std_logic;
          sample_f1_12          : out   std_logic;
          sample_f1_13          : out   std_logic;
          sample_f1_14          : out   std_logic;
          sample_f1_15          : out   std_logic;
          sample_f1_32          : out   std_logic;
          sample_f1_33          : out   std_logic;
          sample_f1_34          : out   std_logic;
          sample_f1_35          : out   std_logic;
          sample_f1_36          : out   std_logic;
          sample_f1_37          : out   std_logic;
          sample_f1_38          : out   std_logic;
          sample_f1_39          : out   std_logic;
          sample_f1_40          : out   std_logic;
          sample_f1_41          : out   std_logic;
          sample_f1_42          : out   std_logic;
          sample_f1_43          : out   std_logic;
          sample_f1_44          : out   std_logic;
          sample_f1_45          : out   std_logic;
          sample_f1_46          : out   std_logic;
          sample_f1_47          : out   std_logic;
          sample_f1_48          : out   std_logic;
          sample_f1_49          : out   std_logic;
          sample_f1_50          : out   std_logic;
          sample_f1_51          : out   std_logic;
          sample_f1_52          : out   std_logic;
          sample_f1_53          : out   std_logic;
          sample_f1_54          : out   std_logic;
          sample_f1_55          : out   std_logic;
          sample_f1_56          : out   std_logic;
          sample_f1_57          : out   std_logic;
          sample_f1_58          : out   std_logic;
          sample_f1_59          : out   std_logic;
          sample_f1_60          : out   std_logic;
          sample_f1_61          : out   std_logic;
          sample_f1_62          : out   std_logic;
          sample_f1_63          : out   std_logic;
          sample_f0_wdata_95    : in    std_logic;
          sample_f0_wdata_94    : in    std_logic;
          sample_f0_wdata_93    : in    std_logic;
          sample_f0_wdata_92    : in    std_logic;
          sample_f0_wdata_91    : in    std_logic;
          sample_f0_wdata_90    : in    std_logic;
          sample_f0_wdata_89    : in    std_logic;
          sample_f0_wdata_88    : in    std_logic;
          sample_f0_wdata_87    : in    std_logic;
          sample_f0_wdata_86    : in    std_logic;
          sample_f0_wdata_85    : in    std_logic;
          sample_f0_wdata_84    : in    std_logic;
          sample_f0_wdata_83    : in    std_logic;
          sample_f0_wdata_82    : in    std_logic;
          sample_f0_wdata_81    : in    std_logic;
          sample_f0_wdata_80    : in    std_logic;
          sample_f0_wdata_79    : in    std_logic;
          sample_f0_wdata_78    : in    std_logic;
          sample_f0_wdata_77    : in    std_logic;
          sample_f0_wdata_76    : in    std_logic;
          sample_f0_wdata_75    : in    std_logic;
          sample_f0_wdata_74    : in    std_logic;
          sample_f0_wdata_73    : in    std_logic;
          sample_f0_wdata_72    : in    std_logic;
          sample_f0_wdata_71    : in    std_logic;
          sample_f0_wdata_70    : in    std_logic;
          sample_f0_wdata_69    : in    std_logic;
          sample_f0_wdata_68    : in    std_logic;
          sample_f0_wdata_67    : in    std_logic;
          sample_f0_wdata_66    : in    std_logic;
          sample_f0_wdata_65    : in    std_logic;
          sample_f0_wdata_64    : in    std_logic;
          sample_f0_wdata_63    : in    std_logic;
          sample_f0_wdata_62    : in    std_logic;
          sample_f0_wdata_61    : in    std_logic;
          sample_f0_wdata_60    : in    std_logic;
          sample_f0_wdata_59    : in    std_logic;
          sample_f0_wdata_58    : in    std_logic;
          sample_f0_wdata_57    : in    std_logic;
          sample_f0_wdata_56    : in    std_logic;
          sample_f0_wdata_55    : in    std_logic;
          sample_f0_wdata_54    : in    std_logic;
          sample_f0_wdata_53    : in    std_logic;
          sample_f0_wdata_52    : in    std_logic;
          sample_f0_wdata_51    : in    std_logic;
          sample_f0_wdata_50    : in    std_logic;
          sample_f0_wdata_49    : in    std_logic;
          sample_f0_wdata_48    : in    std_logic;
          sample_f0_wdata_15    : in    std_logic;
          sample_f0_wdata_14    : in    std_logic;
          sample_f0_wdata_13    : in    std_logic;
          sample_f0_wdata_12    : in    std_logic;
          sample_f0_wdata_11    : in    std_logic;
          sample_f0_wdata_10    : in    std_logic;
          sample_f0_wdata_9     : in    std_logic;
          sample_f0_wdata_8     : in    std_logic;
          sample_f0_wdata_7     : in    std_logic;
          sample_f0_wdata_6     : in    std_logic;
          sample_f0_wdata_5     : in    std_logic;
          sample_f0_wdata_4     : in    std_logic;
          sample_f0_wdata_3     : in    std_logic;
          sample_f0_wdata_2     : in    std_logic;
          sample_f0_wdata_1     : in    std_logic;
          sample_f0_wdata_0     : in    std_logic;
          sample_f1_wdata_95    : out   std_logic;
          sample_f1_wdata_94    : out   std_logic;
          sample_f1_wdata_93    : out   std_logic;
          sample_f1_wdata_92    : out   std_logic;
          sample_f1_wdata_91    : out   std_logic;
          sample_f1_wdata_90    : out   std_logic;
          sample_f1_wdata_89    : out   std_logic;
          sample_f1_wdata_88    : out   std_logic;
          sample_f1_wdata_87    : out   std_logic;
          sample_f1_wdata_86    : out   std_logic;
          sample_f1_wdata_85    : out   std_logic;
          sample_f1_wdata_84    : out   std_logic;
          sample_f1_wdata_83    : out   std_logic;
          sample_f1_wdata_82    : out   std_logic;
          sample_f1_wdata_81    : out   std_logic;
          sample_f1_wdata_80    : out   std_logic;
          sample_f1_wdata_79    : out   std_logic;
          sample_f1_wdata_78    : out   std_logic;
          sample_f1_wdata_77    : out   std_logic;
          sample_f1_wdata_76    : out   std_logic;
          sample_f1_wdata_75    : out   std_logic;
          sample_f1_wdata_74    : out   std_logic;
          sample_f1_wdata_73    : out   std_logic;
          sample_f1_wdata_72    : out   std_logic;
          sample_f1_wdata_71    : out   std_logic;
          sample_f1_wdata_70    : out   std_logic;
          sample_f1_wdata_69    : out   std_logic;
          sample_f1_wdata_68    : out   std_logic;
          sample_f1_wdata_67    : out   std_logic;
          sample_f1_wdata_66    : out   std_logic;
          sample_f1_wdata_65    : out   std_logic;
          sample_f1_wdata_64    : out   std_logic;
          sample_f1_wdata_63    : out   std_logic;
          sample_f1_wdata_62    : out   std_logic;
          sample_f1_wdata_61    : out   std_logic;
          sample_f1_wdata_60    : out   std_logic;
          sample_f1_wdata_59    : out   std_logic;
          sample_f1_wdata_58    : out   std_logic;
          sample_f1_wdata_57    : out   std_logic;
          sample_f1_wdata_56    : out   std_logic;
          sample_f1_wdata_55    : out   std_logic;
          sample_f1_wdata_54    : out   std_logic;
          sample_f1_wdata_53    : out   std_logic;
          sample_f1_wdata_52    : out   std_logic;
          sample_f1_wdata_51    : out   std_logic;
          sample_f1_wdata_50    : out   std_logic;
          sample_f1_wdata_49    : out   std_logic;
          sample_f1_wdata_48    : out   std_logic;
          sample_f1_wdata_15    : out   std_logic;
          sample_f1_wdata_14    : out   std_logic;
          sample_f1_wdata_13    : out   std_logic;
          sample_f1_wdata_12    : out   std_logic;
          sample_f1_wdata_11    : out   std_logic;
          sample_f1_wdata_10    : out   std_logic;
          sample_f1_wdata_9     : out   std_logic;
          sample_f1_wdata_8     : out   std_logic;
          sample_f1_wdata_7     : out   std_logic;
          sample_f1_wdata_6     : out   std_logic;
          sample_f1_wdata_5     : out   std_logic;
          sample_f1_wdata_4     : out   std_logic;
          sample_f1_wdata_3     : out   std_logic;
          sample_f1_wdata_2     : out   std_logic;
          sample_f1_wdata_1     : out   std_logic;
          sample_f1_wdata_0     : out   std_logic;
          sample_f0_val_1       : in    std_logic;
          sample_f1_val         : out   std_logic;
          sample_f0_val_0       : in    std_logic;
          sample_out_0_sqmuxa_1 : out   std_logic;
          HRESETn_c             : in    std_logic;
          HCLK_c                : in    std_logic;
          sample_f1_val_0       : out   std_logic
        );

end Downsampling_8_16_6;

architecture DEF_ARCH of Downsampling_8_16_6 is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal sample_out_val_14, sample_out_0_sqmuxa_3, 
        un10_sample_in_val_24, un10_sample_in_val_25, 
        sample_out_0_sqmuxa_2, sample_out_0_sqmuxa_1_net_1, 
        sample_out_0_sqmuxa_1_0, sample_out_0_sqmuxa_0, 
        un10_sample_in_val_24_0, un10_sample_in_val_15, 
        un10_sample_in_val_14, un10_sample_in_val_20, 
        un10_sample_in_val_25_0, un10_sample_in_val_17, 
        un10_sample_in_val_16, un10_sample_in_val_23, N_137, 
        \counter[1]_net_1\, \counter[0]_net_1\, N_129, 
        \counter[3]_net_1\, \DWACT_FDEC_E[0]\, N_106, 
        \counter[8]_net_1\, \DWACT_FDEC_E[4]\, N_91, 
        \DWACT_FDEC_E[7]\, \DWACT_FDEC_E[6]\, 
        un10_sample_in_val_9, un10_sample_in_val_8, 
        un10_sample_in_val_19, un10_sample_in_val_13, 
        \counter[24]_net_1\, un10_sample_in_val_11, 
        \counter[15]_net_1\, \counter[12]_net_1\, 
        un10_sample_in_val_7, \counter[22]_net_1\, 
        \counter[19]_net_1\, un10_sample_in_val_5, 
        \counter[10]_net_1\, \counter[7]_net_1\, 
        un10_sample_in_val_3, \counter[23]_net_1\, 
        \counter[20]_net_1\, un10_sample_in_val_1, 
        \counter[11]_net_1\, \counter[27]_net_1\, 
        \counter[18]_net_1\, \counter[21]_net_1\, 
        \counter[9]_net_1\, \counter[4]_net_1\, 
        \counter[6]_net_1\, \counter[25]_net_1\, 
        \counter[2]_net_1\, \counter[13]_net_1\, 
        \counter[16]_net_1\, \counter[26]_net_1\, 
        \counter[5]_net_1\, \counter[14]_net_1\, 
        \counter[17]_net_1\, \counter_4[1]\, I_5_0, 
        \counter_4[3]\, I_13_0, \counter_4[4]\, I_20_0, 
        \counter_4[5]\, I_24_0, \counter_4[6]\, I_31_1, 
        \counter_4[7]\, I_38_0, \counter_4[8]\, I_45_0, 
        \counter_4[9]\, I_52_0, \counter_4[10]\, I_56_0, 
        \counter_4[11]\, I_66_0, \counter_4[12]\, I_73_0, 
        \counter_4[13]\, I_77_0, \counter_4[14]\, I_84_0, 
        \counter_4[15]\, I_91_0, \counter_4[16]\, I_98_0, 
        \counter_4[17]\, I_105_0, \counter_4[18]\, I_115_0, 
        \counter_4[19]\, I_122_0, \counter_4[20]\, I_129_0, 
        \counter_4[21]\, I_136_0, \counter_4[22]\, I_143_0, 
        \counter_4[23]\, I_156_0, \counter_4[24]\, I_166_0, 
        \counter_4[25]\, I_173_0, \counter_4[26]\, I_186_0, 
        \counter_4[27]\, I_196_0, sample_out_0_sqmuxa, I_4_0, 
        I_9_0, N_4, \DWACT_FDEC_E[29]\, \DWACT_FDEC_E[30]\, 
        \DWACT_FDEC_E[23]\, \DWACT_FDEC_E[15]\, 
        \DWACT_FDEC_E[17]\, \DWACT_FDEC_E[22]\, N_11, 
        \DWACT_FDEC_E[21]\, \DWACT_FDEC_E[9]\, \DWACT_FDEC_E[12]\, 
        \DWACT_FDEC_E[20]\, N_20, \DWACT_FDEC_E[13]\, 
        \DWACT_FDEC_E[19]\, N_25, \DWACT_FDEC_E[18]\, N_32, 
        \DWACT_FDEC_E[33]\, \DWACT_FDEC_E[34]\, \DWACT_FDEC_E[2]\, 
        \DWACT_FDEC_E[5]\, N_41, \DWACT_FDEC_E[28]\, 
        \DWACT_FDEC_E[16]\, N_46, N_51, \DWACT_FDEC_E[14]\, N_56, 
        N_61, \DWACT_FDEC_E[10]\, N_68, \DWACT_FDEC_E[11]\, N_73, 
        N_78, N_83, \DWACT_FDEC_E[8]\, N_88, N_96, N_103, 
        \DWACT_FDEC_E[3]\, N_111, N_116, N_121, \DWACT_FDEC_E[1]\, 
        N_126, N_134, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    sample_out_0_sqmuxa_1 <= sample_out_0_sqmuxa_1_net_1;

    \counter[19]\ : DFN1E1C0
      port map(D => \counter_4[19]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[19]_net_1\);
    
    \sample_out[125]\ : DFN1E1
      port map(D => sample_f0_wdata_2, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_2);
    
    \sample_out[102]\ : DFN1E1
      port map(D => sample_f0_54, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_54);
    
    \sample_out[122]\ : DFN1E1
      port map(D => sample_f0_wdata_5, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_5);
    
    \sample_out[22]\ : DFN1E1
      port map(D => sample_f0_wdata_73, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_73);
    
    \sample_out[101]\ : DFN1E1
      port map(D => sample_f0_53, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_53);
    
    \sample_out[20]\ : DFN1E1
      port map(D => sample_f0_wdata_75, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_75);
    
    \sample_out[13]\ : DFN1E1
      port map(D => sample_f0_wdata_82, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_82);
    
    \sample_out[1]\ : DFN1E1
      port map(D => sample_f0_wdata_94, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_94);
    
    \sample_out[19]\ : DFN1E1
      port map(D => sample_f0_wdata_76, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_76);
    
    un3_counter_I_142 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[16]\, Y => N_41);
    
    \sample_out[61]\ : DFN1E1
      port map(D => sample_f0_13, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_13);
    
    \sample_out[121]\ : DFN1E1
      port map(D => sample_f0_wdata_6, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_6);
    
    \counter_RNIA89N_0[10]\ : NOR3C
      port map(A => un10_sample_in_val_17, B => 
        un10_sample_in_val_16, C => un10_sample_in_val_23, Y => 
        un10_sample_in_val_25_0);
    
    \sample_out[38]\ : DFN1E1
      port map(D => sample_f0_wdata_57, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_57);
    
    un3_counter_I_27 : OR2
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        Y => \DWACT_FDEC_E[1]\);
    
    \sample_out[95]\ : DFN1E1
      port map(D => sample_f0_47, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_47);
    
    \counter_RNO[11]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_66_0, Y => 
        \counter_4[11]\);
    
    \sample_out[104]\ : DFN1E1
      port map(D => sample_f0_56, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_56);
    
    \sample_out[34]\ : DFN1E1
      port map(D => sample_f0_wdata_61, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_61);
    
    un3_counter_I_4 : INV
      port map(A => \counter[0]_net_1\, Y => I_4_0);
    
    \sample_out[124]\ : DFN1E1
      port map(D => sample_f0_wdata_3, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_3);
    
    \counter[11]\ : DFN1E1C0
      port map(D => \counter_4[11]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[11]_net_1\);
    
    un3_counter_I_94 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, Y
         => \DWACT_FDEC_E[10]\);
    
    \sample_out[97]\ : DFN1E1
      port map(D => sample_f0_49, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_49);
    
    un3_counter_I_186 : XNOR2
      port map(A => N_11, B => \counter[26]_net_1\, Y => I_186_0);
    
    \sample_out[108]\ : DFN1E1
      port map(D => sample_f0_60, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_60);
    
    \counter_RNO[15]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_91_0, Y => \counter_4[15]\);
    
    un3_counter_I_108 : OR3
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        C => \counter[17]_net_1\, Y => \DWACT_FDEC_E[12]\);
    
    un3_counter_I_121 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \counter[18]_net_1\, Y => N_56);
    
    \sample_out[51]\ : DFN1E1
      port map(D => sample_f0_3, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_3);
    
    \sample_out[56]\ : DFN1E1
      port map(D => sample_f0_8, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_8);
    
    un3_counter_I_176 : OR2
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        Y => \DWACT_FDEC_E[20]\);
    
    \sample_out[0]\ : DFN1E1
      port map(D => sample_f0_wdata_95, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_95);
    
    \counter_RNO[7]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_38_0, Y => \counter_4[7]\);
    
    \counter[6]\ : DFN1E1C0
      port map(D => \counter_4[6]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[6]_net_1\);
    
    un3_counter_I_48 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => \DWACT_FDEC_E[4]\);
    
    un3_counter_I_114 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[10]\, 
        C => \DWACT_FDEC_E[12]\, Y => N_61);
    
    \counter[21]\ : DFN1E1C0
      port map(D => \counter_4[21]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[21]_net_1\);
    
    un3_counter_I_13 : XNOR2
      port map(A => N_134, B => \counter[3]_net_1\, Y => I_13_0);
    
    \sample_out[81]\ : DFN1E1
      port map(D => sample_f0_33, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_33);
    
    \sample_out[86]\ : DFN1E1
      port map(D => sample_f0_38, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_38);
    
    \counter[3]\ : DFN1E1C0
      port map(D => \counter_4[3]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[3]_net_1\);
    
    \counter[2]\ : DFN1E1C0
      port map(D => I_9_0, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f0_val_1, Q => \counter[2]_net_1\);
    
    un3_counter_I_73 : XNOR2
      port map(A => N_91, B => \counter[12]_net_1\, Y => I_73_0);
    
    \counter_RNO[8]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_45_0, Y => \counter_4[8]\);
    
    \counter_RNO[13]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_77_0, Y => 
        \counter_4[13]\);
    
    un3_counter_I_52 : XNOR2
      port map(A => N_106, B => \counter[9]_net_1\, Y => I_52_0);
    
    \sample_out[12]\ : DFN1E1
      port map(D => sample_f0_wdata_83, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_83);
    
    \counter_RNINF54[10]\ : NOR3A
      port map(A => un10_sample_in_val_5, B => 
        \counter[10]_net_1\, C => \counter[7]_net_1\, Y => 
        un10_sample_in_val_16);
    
    \sample_out[10]\ : DFN1E1
      port map(D => sample_f0_wdata_85, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_85);
    
    \sample_out[45]\ : DFN1E1
      port map(D => sample_f0_wdata_50, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_50);
    
    \counter_RNO[12]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_73_0, Y => 
        \counter_4[12]\);
    
    \sample_out[33]\ : DFN1E1
      port map(D => sample_f0_wdata_62, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_62);
    
    \sample_out[39]\ : DFN1E1
      port map(D => sample_f0_wdata_56, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_56);
    
    \counter_RNO[1]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_5_0, Y => \counter_4[1]\);
    
    \counter[17]\ : DFN1E1C0
      port map(D => \counter_4[17]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[17]_net_1\);
    
    un3_counter_I_41 : OR2
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        Y => \DWACT_FDEC_E[3]\);
    
    un3_counter_I_159 : OR3
      port map(A => \counter[21]_net_1\, B => \counter[22]_net_1\, 
        C => \counter[23]_net_1\, Y => \DWACT_FDEC_E[17]\);
    
    \counter_RNIRB64[22]\ : NOR3A
      port map(A => un10_sample_in_val_7, B => 
        \counter[22]_net_1\, C => \counter[19]_net_1\, Y => 
        un10_sample_in_val_17);
    
    \counter[4]\ : DFN1E1C0
      port map(D => \counter_4[4]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[4]_net_1\);
    
    un3_counter_I_5 : XNOR2
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        Y => I_5_0);
    
    un3_counter_I_125 : OR2
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        Y => \DWACT_FDEC_E[14]\);
    
    \counter[10]\ : DFN1E1C0
      port map(D => \counter_4[10]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[10]_net_1\);
    
    \sample_out[5]\ : DFN1E1
      port map(D => sample_f0_wdata_90, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_wdata_90);
    
    \sample_out[47]\ : DFN1E1
      port map(D => sample_f0_wdata_48, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_wdata_48);
    
    \counter_RNI91T[12]\ : NOR3A
      port map(A => un10_sample_in_val_11, B => 
        \counter[15]_net_1\, C => \counter[12]_net_1\, Y => 
        un10_sample_in_val_19);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter[13]\ : DFN1E1C0
      port map(D => \counter_4[13]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[13]_net_1\);
    
    un3_counter_I_62 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[6]\);
    
    un3_counter_I_139 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        Y => \DWACT_FDEC_E[16]\);
    
    \sample_out[115]\ : DFN1E1
      port map(D => sample_f0_wdata_12, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_12);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sample_out[21]\ : DFN1E1
      port map(D => sample_f0_wdata_74, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_74);
    
    \counter[12]\ : DFN1E1C0
      port map(D => \counter_4[12]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[12]_net_1\);
    
    \sample_out[26]\ : DFN1E1
      port map(D => sample_f0_wdata_69, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_69);
    
    \sample_out[2]\ : DFN1E1
      port map(D => sample_f0_wdata_93, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_93);
    
    \sample_out[98]\ : DFN1E1
      port map(D => sample_f0_50, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_50);
    
    \sample_out[112]\ : DFN1E1
      port map(D => sample_f0_wdata_15, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_15);
    
    \counter[27]\ : DFN1E1C0
      port map(D => \counter_4[27]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[27]_net_1\);
    
    \counter_RNIIDQF[20]\ : NOR3C
      port map(A => un10_sample_in_val_15, B => 
        un10_sample_in_val_14, C => un10_sample_in_val_20, Y => 
        un10_sample_in_val_24);
    
    un3_counter_I_111 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[28]\);
    
    \counter[20]\ : DFN1E1C0
      port map(D => \counter_4[20]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[20]_net_1\);
    
    \sample_out[94]\ : DFN1E1
      port map(D => sample_f0_46, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_46);
    
    \sample_out[111]\ : DFN1E1
      port map(D => sample_f0_63, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_63);
    
    \counter_RNIMKE[21]\ : NOR2
      port map(A => \counter[18]_net_1\, B => \counter[21]_net_1\, 
        Y => un10_sample_in_val_11);
    
    un3_counter_I_166 : XNOR2
      port map(A => N_25, B => \counter[24]_net_1\, Y => I_166_0);
    
    \counter_RNO[17]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_105_0, Y => \counter_4[17]\);
    
    \counter[23]\ : DFN1E1C0
      port map(D => \counter_4[23]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[23]_net_1\);
    
    un3_counter_I_149 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[34]\);
    
    \sample_out[55]\ : DFN1E1
      port map(D => sample_f0_7, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_7);
    
    \counter[22]\ : DFN1E1C0
      port map(D => \counter_4[22]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[22]_net_1\);
    
    \counter[15]\ : DFN1E1C0
      port map(D => \counter_4[15]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[15]_net_1\);
    
    un3_counter_I_8 : OR2
      port map(A => \counter[1]_net_1\, B => \counter[0]_net_1\, 
        Y => N_137);
    
    un3_counter_I_185 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[21]\, Y => N_11);
    
    \sample_out[114]\ : DFN1E1
      port map(D => sample_f0_wdata_13, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_13);
    
    un3_counter_I_196 : XNOR2
      port map(A => N_4, B => \counter[27]_net_1\, Y => I_196_0);
    
    \sample_out[32]\ : DFN1E1
      port map(D => sample_f0_wdata_63, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_63);
    
    un3_counter_I_51 : OR2
      port map(A => \counter[8]_net_1\, B => \DWACT_FDEC_E[4]\, Y
         => N_106);
    
    un3_counter_I_122 : XNOR2
      port map(A => N_56, B => \counter[19]_net_1\, Y => I_122_0);
    
    \counter_RNILKE[13]\ : NOR2
      port map(A => \counter[13]_net_1\, B => \counter[16]_net_1\, 
        Y => un10_sample_in_val_5);
    
    \sample_out[118]\ : DFN1E1
      port map(D => sample_f0_wdata_9, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_9);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sample_out[57]\ : DFN1E1
      port map(D => sample_f0_9, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_9);
    
    \sample_out[30]\ : DFN1E1
      port map(D => sample_f0_wdata_65, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_65);
    
    \counter_RNO[14]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_84_0, Y => 
        \counter_4[14]\);
    
    \sample_out[85]\ : DFN1E1
      port map(D => sample_f0_37, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_37);
    
    \counter[1]\ : DFN1E1C0
      port map(D => \counter_4[1]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[1]_net_1\);
    
    \counter_RNO[26]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_186_0, Y => \counter_4[26]\);
    
    \sample_out[4]\ : DFN1E1
      port map(D => sample_f0_wdata_91, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_wdata_91);
    
    \counter_RNO[5]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_24_0, Y => \counter_4[5]\);
    
    \sample_out[103]\ : DFN1E1
      port map(D => sample_f0_55, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_55);
    
    \sample_out[100]\ : DFN1E1
      port map(D => sample_f0_52, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_52);
    
    \counter_RNI7KBF1_0[10]\ : NOR3C
      port map(A => un10_sample_in_val_24, B => 
        un10_sample_in_val_25, C => sample_out_0_sqmuxa_1_net_1, 
        Y => sample_out_0_sqmuxa_2);
    
    \counter[25]\ : DFN1E1C0
      port map(D => \counter_4[25]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[25]_net_1\);
    
    \sample_out[123]\ : DFN1E1
      port map(D => sample_f0_wdata_4, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_4);
    
    \sample_out[120]\ : DFN1E1
      port map(D => sample_f0_wdata_7, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_7);
    
    sample_out_val : DFN1C0
      port map(D => sample_out_val_14, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f1_val);
    
    \counter_RNO[3]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_13_0, Y => \counter_4[3]\);
    
    \sample_out[87]\ : DFN1E1
      port map(D => sample_f0_39, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_39);
    
    un3_counter_I_115 : XNOR2
      port map(A => N_61, B => \counter[18]_net_1\, Y => I_115_0);
    
    un3_counter_I_87 : OR3
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        C => \counter[14]_net_1\, Y => \DWACT_FDEC_E[9]\);
    
    un3_counter_I_173 : XNOR2
      port map(A => N_20, B => \counter[25]_net_1\, Y => I_173_0);
    
    \sample_out[48]\ : DFN1E1
      port map(D => sample_f0_0, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_0);
    
    un3_counter_I_38 : XNOR2
      port map(A => N_116, B => \counter[7]_net_1\, Y => I_38_0);
    
    \counter_RNID507[3]\ : NOR2
      port map(A => \counter[3]_net_1\, B => \counter[0]_net_1\, 
        Y => un10_sample_in_val_13);
    
    \sample_out[93]\ : DFN1E1
      port map(D => sample_f0_45, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_45);
    
    \sample_out[11]\ : DFN1E1
      port map(D => sample_f0_wdata_84, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_84);
    
    \sample_out[99]\ : DFN1E1
      port map(D => sample_f0_51, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_51);
    
    \sample_out[16]\ : DFN1E1
      port map(D => sample_f0_wdata_79, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_79);
    
    \counter[5]\ : DFN1E1C0
      port map(D => \counter_4[5]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[5]_net_1\);
    
    \sample_out[44]\ : DFN1E1
      port map(D => sample_f0_wdata_51, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_51);
    
    un3_counter_I_37 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \counter[6]_net_1\, Y => N_116);
    
    \counter_RNO[10]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_56_0, Y => 
        \counter_4[10]\);
    
    un3_counter_I_9 : XNOR2
      port map(A => N_137, B => \counter[2]_net_1\, Y => I_9_0);
    
    \counter_RNO[21]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_136_0, Y => \counter_4[21]\);
    
    un3_counter_I_20 : XNOR2
      port map(A => N_129, B => \counter[4]_net_1\, Y => I_20_0);
    
    \counter_RNIK507[4]\ : NOR2
      port map(A => \counter[4]_net_1\, B => \counter[6]_net_1\, 
        Y => un10_sample_in_val_8);
    
    un3_counter_I_182 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[30]\);
    
    \sample_out[25]\ : DFN1E1
      port map(D => sample_f0_wdata_70, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_70);
    
    \counter_RNI7KBF1_3[10]\ : NOR3C
      port map(A => un10_sample_in_val_24, B => 
        un10_sample_in_val_25, C => sample_out_0_sqmuxa_1_net_1, 
        Y => sample_out_0_sqmuxa);
    
    un3_counter_I_56 : XNOR2
      port map(A => N_103, B => \counter[10]_net_1\, Y => I_56_0);
    
    \counter[16]\ : DFN1E1C0
      port map(D => \counter_4[16]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[16]_net_1\);
    
    \counter_RNO[25]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_173_0, Y => \counter_4[25]\);
    
    un3_counter_I_172 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[19]\, Y => N_20);
    
    un3_counter_I_104 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \DWACT_FDEC_E[11]\, Y => N_68);
    
    un3_counter_I_31 : XNOR2
      port map(A => N_121, B => \counter[6]_net_1\, Y => I_31_1);
    
    un3_counter_I_98 : XNOR2
      port map(A => N_73, B => \counter[16]_net_1\, Y => I_98_0);
    
    un3_counter_I_23 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \counter[3]_net_1\, C
         => \counter[4]_net_1\, Y => N_126);
    
    \sample_out[27]\ : DFN1E1
      port map(D => sample_f0_wdata_68, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_68);
    
    un3_counter_I_59 : OR3
      port map(A => \counter[6]_net_1\, B => \counter[7]_net_1\, 
        C => \counter[8]_net_1\, Y => \DWACT_FDEC_E[5]\);
    
    un3_counter_I_12 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => N_134);
    
    \counter_RNO[6]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_31_1, Y => \counter_4[6]\);
    
    un3_counter_I_165 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[18]\, Y => N_25);
    
    un3_counter_I_156 : XNOR2
      port map(A => N_32, B => \counter[23]_net_1\, Y => I_156_0);
    
    un3_counter_I_97 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[10]\, C
         => \counter[15]_net_1\, Y => N_73);
    
    un3_counter_I_128 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[14]\, Y => N_51);
    
    un3_counter_I_72 : OR2
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[6]\, Y
         => N_91);
    
    \sample_out[58]\ : DFN1E1
      port map(D => sample_f0_10, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_10);
    
    \counter[26]\ : DFN1E1C0
      port map(D => \counter_4[26]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[26]_net_1\);
    
    un3_counter_I_66 : XNOR2
      port map(A => N_96, B => \counter[11]_net_1\, Y => I_66_0);
    
    \counter_RNO[23]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_156_0, Y => \counter_4[23]\);
    
    \sample_out[54]\ : DFN1E1
      port map(D => sample_f0_6, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_6);
    
    \sample_out[43]\ : DFN1E1
      port map(D => sample_f0_wdata_52, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_52);
    
    \sample_out[49]\ : DFN1E1
      port map(D => sample_f0_1, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_1);
    
    sample_out_val_0 : DFN1C0
      port map(D => sample_out_val_14, CLK => HCLK_c, CLR => 
        HRESETn_c, Q => sample_f1_val_0);
    
    \counter_RNI3FN3[25]\ : NOR2
      port map(A => \counter[25]_net_1\, B => \counter[2]_net_1\, 
        Y => un10_sample_in_val_7);
    
    un3_counter_I_45 : XNOR2
      port map(A => N_111, B => \counter[8]_net_1\, Y => I_45_0);
    
    un3_counter_I_24 : XNOR2
      port map(A => N_126, B => \counter[5]_net_1\, Y => I_24_0);
    
    un3_counter_I_195 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[30]\, 
        C => \DWACT_FDEC_E[23]\, Y => N_4);
    
    \sample_out[92]\ : DFN1E1
      port map(D => sample_f0_44, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_44);
    
    \counter[14]\ : DFN1E1C0
      port map(D => \counter_4[14]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[14]_net_1\);
    
    un3_counter_I_136 : XNOR2
      port map(A => N_46, B => \counter[21]_net_1\, Y => I_136_0);
    
    \sample_out[88]\ : DFN1E1
      port map(D => sample_f0_40, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_40);
    
    \sample_out[90]\ : DFN1E1
      port map(D => sample_f0_42, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_42);
    
    un3_counter_I_91 : XNOR2
      port map(A => N_78, B => \counter[15]_net_1\, Y => I_91_0);
    
    \counter_RNO[22]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_143_0, Y => \counter_4[22]\);
    
    \sample_out[31]\ : DFN1E1
      port map(D => sample_f0_wdata_64, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_64);
    
    \sample_out[36]\ : DFN1E1
      port map(D => sample_f0_wdata_59, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_59);
    
    un3_counter_I_69 : OR3
      port map(A => \counter[9]_net_1\, B => \counter[10]_net_1\, 
        C => \counter[11]_net_1\, Y => \DWACT_FDEC_E[7]\);
    
    \sample_out_0_sqmuxa_1\ : NOR2B
      port map(A => sample_f0_val_0, B => HRESETn_c, Y => 
        sample_out_0_sqmuxa_1_net_1);
    
    \sample_out[84]\ : DFN1E1
      port map(D => sample_f0_36, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_36);
    
    \sample_out[63]\ : DFN1E1
      port map(D => sample_f0_15, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_15);
    
    \sample_out[15]\ : DFN1E1
      port map(D => sample_f0_wdata_80, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_80);
    
    un3_counter_I_129 : XNOR2
      port map(A => N_51, B => \counter[20]_net_1\, Y => I_129_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    un3_counter_I_146 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \counter[21]_net_1\, 
        C => \counter[22]_net_1\, Y => \DWACT_FDEC_E[33]\);
    
    \counter[24]\ : DFN1E1C0
      port map(D => \counter_4[24]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[24]_net_1\);
    
    un3_counter_I_101 : OR2
      port map(A => \counter[15]_net_1\, B => \counter[16]_net_1\, 
        Y => \DWACT_FDEC_E[11]\);
    
    \sample_out[113]\ : DFN1E1
      port map(D => sample_f0_wdata_14, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_14);
    
    \sample_out[110]\ : DFN1E1
      port map(D => sample_f0_62, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_62);
    
    \counter_RNO[4]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_20_0, Y => \counter_4[4]\);
    
    un3_counter_I_162 : OR2
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        Y => \DWACT_FDEC_E[18]\);
    
    \counter_RNI7KBF1_1[10]\ : NOR3C
      port map(A => un10_sample_in_val_24, B => 
        un10_sample_in_val_25, C => sample_out_0_sqmuxa_1_net_1, 
        Y => sample_out_0_sqmuxa_0);
    
    \counter_RNINSE[14]\ : NOR2
      port map(A => \counter[14]_net_1\, B => \counter[17]_net_1\, 
        Y => un10_sample_in_val_1);
    
    \sample_out[106]\ : DFN1E1
      port map(D => sample_f0_58, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_58);
    
    un3_counter_I_77 : XNOR2
      port map(A => N_88, B => \counter[13]_net_1\, Y => I_77_0);
    
    \sample_out[17]\ : DFN1E1
      port map(D => sample_f0_wdata_78, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_78);
    
    \sample_out[107]\ : DFN1E1
      port map(D => sample_f0_59, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_59);
    
    \counter_RNO[18]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_115_0, Y => \counter_4[18]\);
    
    un3_counter_I_44 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[3]\, Y => N_111);
    
    \sample_out[126]\ : DFN1E1
      port map(D => sample_f0_wdata_1, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_1);
    
    \sample_out[127]\ : DFN1E1
      port map(D => sample_f0_wdata_0, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_0);
    
    \sample_out[53]\ : DFN1E1
      port map(D => sample_f0_5, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_5);
    
    \sample_out[28]\ : DFN1E1
      port map(D => sample_f0_wdata_67, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_67);
    
    \counter_RNO[27]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_196_0, Y => \counter_4[27]\);
    
    \sample_out[59]\ : DFN1E1
      port map(D => sample_f0_11, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_11);
    
    \counter_RNI7KBF1_2[10]\ : NOR3C
      port map(A => un10_sample_in_val_24, B => 
        un10_sample_in_val_25, C => sample_out_0_sqmuxa_1_net_1, 
        Y => sample_out_0_sqmuxa_3);
    
    \sample_out[109]\ : DFN1E1
      port map(D => sample_f0_61, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_61);
    
    un3_counter_I_192 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[22]\, Y => \DWACT_FDEC_E[23]\);
    
    \sample_out[24]\ : DFN1E1
      port map(D => sample_f0_wdata_71, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_71);
    
    \counter_RNIOF54[20]\ : NOR3A
      port map(A => un10_sample_in_val_3, B => 
        \counter[23]_net_1\, C => \counter[20]_net_1\, Y => 
        un10_sample_in_val_15);
    
    \counter_RNIOCTE[12]\ : NOR3C
      port map(A => un10_sample_in_val_9, B => 
        un10_sample_in_val_8, C => un10_sample_in_val_19, Y => 
        un10_sample_in_val_23);
    
    un3_counter_I_55 : OR3
      port map(A => \DWACT_FDEC_E[4]\, B => \counter[8]_net_1\, C
         => \counter[9]_net_1\, Y => N_103);
    
    \sample_out[42]\ : DFN1E1
      port map(D => sample_f0_wdata_53, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_53);
    
    un3_counter_I_118 : OR3
      port map(A => \DWACT_FDEC_E[7]\, B => \DWACT_FDEC_E[9]\, C
         => \DWACT_FDEC_E[12]\, Y => \DWACT_FDEC_E[13]\);
    
    \sample_out[40]\ : DFN1E1
      port map(D => sample_f0_wdata_55, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_55);
    
    \sample_out[83]\ : DFN1E1
      port map(D => sample_f0_35, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_35);
    
    \sample_out[89]\ : DFN1E1
      port map(D => sample_f0_41, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_41);
    
    un3_counter_I_189 : OR3
      port map(A => \counter[24]_net_1\, B => \counter[25]_net_1\, 
        C => \counter[26]_net_1\, Y => \DWACT_FDEC_E[22]\);
    
    \counter_RNO[24]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_166_0, Y => \counter_4[24]\);
    
    \counter[7]\ : DFN1E1C0
      port map(D => \counter_4[7]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[7]_net_1\);
    
    un3_counter_I_105 : XNOR2
      port map(A => N_68, B => \counter[17]_net_1\, Y => I_105_0);
    
    \sample_out[6]\ : DFN1E1
      port map(D => sample_f0_wdata_89, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_wdata_89);
    
    un3_counter_I_155 : OR3
      port map(A => \DWACT_FDEC_E[29]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[33]\, Y => N_32);
    
    un3_counter_I_179 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \DWACT_FDEC_E[20]\, Y => \DWACT_FDEC_E[21]\);
    
    \sample_out[62]\ : DFN1E1
      port map(D => sample_f0_14, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_14);
    
    \sample_out[60]\ : DFN1E1
      port map(D => sample_f0_12, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_12);
    
    un3_counter_I_65 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \counter[9]_net_1\, C
         => \counter[10]_net_1\, Y => N_96);
    
    \counter_RNI7JN3[26]\ : NOR2
      port map(A => \counter[26]_net_1\, B => \counter[5]_net_1\, 
        Y => un10_sample_in_val_3);
    
    \sample_out[35]\ : DFN1E1
      port map(D => sample_f0_wdata_60, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_60);
    
    \sample_out[91]\ : DFN1E1
      port map(D => sample_f0_43, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_43);
    
    un3_counter_I_135 : OR3
      port map(A => \DWACT_FDEC_E[28]\, B => \DWACT_FDEC_E[13]\, 
        C => \DWACT_FDEC_E[15]\, Y => N_46);
    
    \sample_out[96]\ : DFN1E1
      port map(D => sample_f0_48, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_48);
    
    \counter_RNICDT[27]\ : NOR3A
      port map(A => un10_sample_in_val_1, B => 
        \counter[11]_net_1\, C => \counter[27]_net_1\, Y => 
        un10_sample_in_val_14);
    
    un3_counter_I_80 : OR2
      port map(A => \counter[12]_net_1\, B => \counter[13]_net_1\, 
        Y => \DWACT_FDEC_E[8]\);
    
    \counter_RNI8A2C1[10]\ : NOR3C
      port map(A => un10_sample_in_val_24_0, B => 
        un10_sample_in_val_25_0, C => sample_f0_val_0, Y => 
        sample_out_val_14);
    
    un3_counter_I_16 : OR3
      port map(A => \counter[0]_net_1\, B => \counter[1]_net_1\, 
        C => \counter[2]_net_1\, Y => \DWACT_FDEC_E[0]\);
    
    \counter_RNO[20]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_129_0, Y => \counter_4[20]\);
    
    \sample_out[37]\ : DFN1E1
      port map(D => sample_f0_wdata_58, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_58);
    
    \sample_out[23]\ : DFN1E1
      port map(D => sample_f0_wdata_72, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_72);
    
    \sample_out[52]\ : DFN1E1
      port map(D => sample_f0_4, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_4);
    
    \sample_out[29]\ : DFN1E1
      port map(D => sample_f0_wdata_66, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_66);
    
    \counter_RNIEGNA[24]\ : NOR3A
      port map(A => un10_sample_in_val_13, B => 
        \counter[1]_net_1\, C => \counter[24]_net_1\, Y => 
        un10_sample_in_val_20);
    
    un3_counter_I_76 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \counter[12]_net_1\, Y => N_88);
    
    un3_counter_I_30 : OR3
      port map(A => \DWACT_FDEC_E[0]\, B => \DWACT_FDEC_E[1]\, C
         => \counter[5]_net_1\, Y => N_121);
    
    \sample_out[50]\ : DFN1E1
      port map(D => sample_f0_2, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_2);
    
    \sample_out[18]\ : DFN1E1
      port map(D => sample_f0_wdata_77, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_77);
    
    \sample_out[9]\ : DFN1E1
      port map(D => sample_f0_wdata_86, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_wdata_86);
    
    \sample_out[7]\ : DFN1E1
      port map(D => sample_f0_wdata_88, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_wdata_88);
    
    un3_counter_I_83 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[8]\, Y => N_83);
    
    un3_counter_I_19 : OR2
      port map(A => \counter[3]_net_1\, B => \DWACT_FDEC_E[0]\, Y
         => N_129);
    
    \sample_out[14]\ : DFN1E1
      port map(D => sample_f0_wdata_81, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_1_0, Q => sample_f1_wdata_81);
    
    \counter_RNI7KBF1[10]\ : NOR3C
      port map(A => un10_sample_in_val_24, B => 
        un10_sample_in_val_25, C => sample_out_0_sqmuxa_1_net_1, 
        Y => sample_out_0_sqmuxa_1_0);
    
    \sample_out[82]\ : DFN1E1
      port map(D => sample_f0_34, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_34);
    
    \counter[9]\ : DFN1E1C0
      port map(D => \counter_4[9]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[9]_net_1\);
    
    \counter_RNIA89N[10]\ : NOR3C
      port map(A => un10_sample_in_val_17, B => 
        un10_sample_in_val_16, C => un10_sample_in_val_23, Y => 
        un10_sample_in_val_25);
    
    \sample_out[80]\ : DFN1E1
      port map(D => sample_f0_32, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_3, Q => sample_f1_32);
    
    \counter_RNO[19]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_122_0, Y => \counter_4[19]\);
    
    un3_counter_I_152 : OR3
      port map(A => \DWACT_FDEC_E[34]\, B => \DWACT_FDEC_E[2]\, C
         => \DWACT_FDEC_E[5]\, Y => \DWACT_FDEC_E[29]\);
    
    \counter_RNO[9]\ : AOI1B
      port map(A => un10_sample_in_val_25_0, B => 
        un10_sample_in_val_24_0, C => I_52_0, Y => \counter_4[9]\);
    
    \counter[8]\ : DFN1E1C0
      port map(D => \counter_4[8]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_1, Q => \counter[8]_net_1\);
    
    un3_counter_I_84 : XNOR2
      port map(A => N_83, B => \counter[14]_net_1\, Y => I_84_0);
    
    un3_counter_I_143 : XNOR2
      port map(A => N_41, B => \counter[22]_net_1\, Y => I_143_0);
    
    \counter_RNIR507[8]\ : NOR2
      port map(A => \counter[8]_net_1\, B => \counter[9]_net_1\, 
        Y => un10_sample_in_val_9);
    
    \sample_out[116]\ : DFN1E1
      port map(D => sample_f0_wdata_11, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_11);
    
    \counter[18]\ : DFN1E1C0
      port map(D => \counter_4[18]\, CLK => HCLK_c, CLR => 
        HRESETn_c, E => sample_f0_val_0, Q => \counter[18]_net_1\);
    
    \sample_out[117]\ : DFN1E1
      port map(D => sample_f0_wdata_10, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_10);
    
    un3_counter_I_90 : OR3
      port map(A => \DWACT_FDEC_E[6]\, B => \DWACT_FDEC_E[7]\, C
         => \DWACT_FDEC_E[9]\, Y => N_78);
    
    un3_counter_I_169 : OR3
      port map(A => \DWACT_FDEC_E[15]\, B => \DWACT_FDEC_E[17]\, 
        C => \counter[24]_net_1\, Y => \DWACT_FDEC_E[19]\);
    
    un3_counter_I_132 : OR3
      port map(A => \counter[18]_net_1\, B => \counter[19]_net_1\, 
        C => \counter[20]_net_1\, Y => \DWACT_FDEC_E[15]\);
    
    \counter_RNIIDQF_0[20]\ : NOR3C
      port map(A => un10_sample_in_val_15, B => 
        un10_sample_in_val_14, C => un10_sample_in_val_20, Y => 
        un10_sample_in_val_24_0);
    
    \sample_out[8]\ : DFN1E1
      port map(D => sample_f0_wdata_87, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa, Q => sample_f1_wdata_87);
    
    \sample_out[41]\ : DFN1E1
      port map(D => sample_f0_wdata_54, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_54);
    
    \counter_RNO[16]\ : AOI1B
      port map(A => un10_sample_in_val_25, B => 
        un10_sample_in_val_24, C => I_98_0, Y => \counter_4[16]\);
    
    \counter[0]\ : DFN1E1C0
      port map(D => I_4_0, CLK => HCLK_c, CLR => HRESETn_c, E => 
        sample_f0_val_0, Q => \counter[0]_net_1\);
    
    \sample_out[46]\ : DFN1E1
      port map(D => sample_f0_wdata_49, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_49);
    
    \sample_out[3]\ : DFN1E1
      port map(D => sample_f0_wdata_92, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_2, Q => sample_f1_wdata_92);
    
    un3_counter_I_34 : OR3
      port map(A => \counter[3]_net_1\, B => \counter[4]_net_1\, 
        C => \counter[5]_net_1\, Y => \DWACT_FDEC_E[2]\);
    
    \sample_out[105]\ : DFN1E1
      port map(D => sample_f0_57, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_57);
    
    \sample_out[119]\ : DFN1E1
      port map(D => sample_f0_wdata_8, CLK => HCLK_c, E => 
        sample_out_0_sqmuxa_0, Q => sample_f1_wdata_8);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_FF_1 is

    port( cnv_run_c    : in    std_logic;
          HRESETn_c    : in    std_logic;
          HCLK_c       : in    std_logic;
          cnv_run_sync : out   std_logic
        );

end SYNC_FF_1;

architecture DEF_ARCH of SYNC_FF_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \A_temp[1]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sync_loop.0.A_temp[0]\ : DFN1C0
      port map(D => \A_temp[1]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => cnv_run_sync);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \sync_loop.1.A_temp[1]\ : DFN1C0
      port map(D => cnv_run_c, CLK => HCLK_c, CLR => HRESETn_c, Q
         => \A_temp[1]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_FF is

    port( cnv_c      : in    std_logic;
          HRESETn_c  : in    std_logic;
          HCLK_c     : in    std_logic;
          cnv_sync   : out   std_logic;
          cnv_sync_i : out   std_logic
        );

end SYNC_FF;

architecture DEF_ARCH of SYNC_FF is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \cnv_sync\, \A_temp[1]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    cnv_sync <= \cnv_sync\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \sync_loop.0.A_temp[0]\ : DFN1C0
      port map(D => \A_temp[1]\, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => \cnv_sync\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \sync_loop.1.A_temp[1]\ : DFN1C0
      port map(D => cnv_c, CLK => HCLK_c, CLR => HRESETn_c, Q => 
        \A_temp[1]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sync_loop.0.A_temp_RNIEBA5[0]\ : INV
      port map(A => \cnv_sync\, Y => cnv_sync_i);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity AD7688_drvr is

    port( sample_7   : out   std_logic_vector(15 downto 0);
          sample_0   : out   std_logic_vector(15 downto 0);
          sample_1   : out   std_logic_vector(15 downto 0);
          sample_2   : out   std_logic_vector(15 downto 0);
          sample_3   : out   std_logic_vector(15 downto 0);
          sample_4   : out   std_logic_vector(15 downto 0);
          sample_5   : out   std_logic_vector(15 downto 0);
          sdo_c      : in    std_logic_vector(7 downto 0);
          sample_6   : out   std_logic_vector(15 downto 0);
          cnv_rstn_c : in    std_logic;
          cnv_clk_c  : in    std_logic;
          cnv_c      : out   std_logic;
          sample_val : out   std_logic;
          sck_c      : out   std_logic;
          cnv_run_c  : in    std_logic;
          HRESETn_c  : in    std_logic;
          HCLK_c     : in    std_logic
        );

end AD7688_drvr;

architecture DEF_ARCH of AD7688_drvr is 

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SYNC_FF_1
    port( cnv_run_c    : in    std_logic := 'U';
          HRESETn_c    : in    std_logic := 'U';
          HCLK_c       : in    std_logic := 'U';
          cnv_run_sync : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SYNC_FF
    port( cnv_c      : in    std_logic := 'U';
          HRESETn_c  : in    std_logic := 'U';
          HCLK_c     : in    std_logic := 'U';
          cnv_sync   : out   std_logic;
          cnv_sync_i : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sample_bit_counter_4[0]_net_1\, 
        sample_bit_counter_n0, N_6, 
        \sample_bit_counter_3[0]_net_1\, 
        \sample_bit_counter_2[0]_net_1\, 
        \sample_bit_counter_1[0]_net_1\, 
        \sample_bit_counter_0[0]_net_1\, sample_0_0_sqmuxa, 
        \sample_bit_counter_RNIVMI9[5]_net_1\, 
        \sample_bit_counter_i[0]\, sample_bit_counterlde_i_a3_0_1, 
        \sample_bit_counter[3]_net_1\, 
        \sample_bit_counter[2]_net_1\, 
        \sample_bit_counter[4]_net_1\, un3_cnv_runlto8_0, 
        \cnv_cycle_counter[8]_net_1\, 
        \cnv_cycle_counter[7]_net_1\, un3_cnv_runlto5_0, 
        \cnv_cycle_counter[4]_net_1\, 
        \cnv_cycle_counter[5]_net_1\, un2_cnv_runlto8_2, 
        \cnv_cycle_counter[2]_net_1\, 
        \cnv_cycle_counter[3]_net_1\, un2_cnv_runlto8_1, 
        \cnv_cycle_counter[6]_net_1\, un2_cnv_runlto8_0, N_30, 
        N_38, N_36, N_17, N_22, N_15, N_21, N_13, N_20, N_11, 
        un3_cnv_runlt6, cnv_cycle_counter_c2, un3_cnv_run, 
        un2_cnv_run, cnv_cycle_counter_n8, cnv_cycle_counter_33_0, 
        cnv_s_0_sqmuxa, cnv_cycle_counter_n7, 
        cnv_cycle_counter_c6, cnv_cycle_counter_n6, 
        cnv_cycle_counter_c5, cnv_cycle_counter_n5, 
        cnv_cycle_counter_c4, cnv_cycle_counter_n4, 
        cnv_cycle_counter_n4_tz_i, cnv_cycle_counter_n3, 
        cnv_cycle_counter_n3_tz_i, cnv_cycle_counter_n2, 
        cnv_cycle_counter_n2_tz_i, \cnv_cycle_counter[0]_net_1\, 
        \cnv_cycle_counter[1]_net_1\, N_23, 
        \sample_bit_counter[1]_net_1\, N_19, cnv_done_i, 
        cnv_run_sync, \sample_bit_counter[5]_net_1\, 
        \sample_bit_counter_RNI0D96[5]_net_1\, 
        cnv_cycle_counter_n1, cnv_cycle_counter_n0, \cnv_s_RNO\, 
        cnv_done_1, cnv_sync_r_i_0, cnv_sync, cnv_sync_i, 
        \sample_bit_counter[0]_net_1\, \shift_reg_6[0]_net_1\, 
        \shift_reg_6[1]_net_1\, \shift_reg_6[2]_net_1\, 
        \shift_reg_6[3]_net_1\, \shift_reg_6[4]_net_1\, 
        \shift_reg_6[5]_net_1\, \shift_reg_6[6]_net_1\, 
        \shift_reg_6[7]_net_1\, \shift_reg_6[8]_net_1\, 
        \shift_reg_6[9]_net_1\, \shift_reg_6[10]_net_1\, 
        \shift_reg_6[11]_net_1\, \shift_reg_6[12]_net_1\, 
        \shift_reg_6[13]_net_1\, \shift_reg_6[14]_net_1\, 
        \shift_reg_5[0]_net_1\, \shift_reg_5[1]_net_1\, 
        \shift_reg_5[2]_net_1\, \shift_reg_5[3]_net_1\, 
        \shift_reg_5[4]_net_1\, \shift_reg_5[5]_net_1\, 
        \shift_reg_5[6]_net_1\, \shift_reg_5[7]_net_1\, 
        \shift_reg_5[8]_net_1\, \shift_reg_5[9]_net_1\, 
        \shift_reg_5[10]_net_1\, \shift_reg_5[11]_net_1\, 
        \shift_reg_5[12]_net_1\, \shift_reg_5[13]_net_1\, 
        \shift_reg_5[14]_net_1\, \shift_reg_4[0]_net_1\, 
        \shift_reg_4[1]_net_1\, \shift_reg_4[2]_net_1\, 
        \shift_reg_4[3]_net_1\, \shift_reg_4[4]_net_1\, 
        \shift_reg_4[5]_net_1\, \shift_reg_4[6]_net_1\, 
        \shift_reg_4[7]_net_1\, \shift_reg_4[8]_net_1\, 
        \shift_reg_4[9]_net_1\, \shift_reg_4[10]_net_1\, 
        \shift_reg_4[11]_net_1\, \shift_reg_4[12]_net_1\, 
        \shift_reg_4[13]_net_1\, \shift_reg_4[14]_net_1\, 
        \shift_reg_3[0]_net_1\, \shift_reg_3[1]_net_1\, 
        \shift_reg_3[2]_net_1\, \shift_reg_3[3]_net_1\, 
        \shift_reg_3[4]_net_1\, \shift_reg_3[5]_net_1\, 
        \shift_reg_3[6]_net_1\, \shift_reg_3[7]_net_1\, 
        \shift_reg_3[8]_net_1\, \shift_reg_3[9]_net_1\, 
        \shift_reg_3[10]_net_1\, \shift_reg_3[11]_net_1\, 
        \shift_reg_3[12]_net_1\, \shift_reg_3[13]_net_1\, 
        \shift_reg_3[14]_net_1\, \shift_reg_2[0]_net_1\, 
        \shift_reg_2[1]_net_1\, \shift_reg_2[2]_net_1\, 
        \shift_reg_2[3]_net_1\, \shift_reg_2[4]_net_1\, 
        \shift_reg_2[5]_net_1\, \shift_reg_2[6]_net_1\, 
        \shift_reg_2[7]_net_1\, \shift_reg_2[8]_net_1\, 
        \shift_reg_2[9]_net_1\, \shift_reg_2[10]_net_1\, 
        \shift_reg_2[11]_net_1\, \shift_reg_2[12]_net_1\, 
        \shift_reg_2[13]_net_1\, \shift_reg_2[14]_net_1\, 
        \shift_reg_1[0]_net_1\, \shift_reg_1[1]_net_1\, 
        \shift_reg_1[2]_net_1\, \shift_reg_1[3]_net_1\, 
        \shift_reg_1[4]_net_1\, \shift_reg_1[5]_net_1\, 
        \shift_reg_1[6]_net_1\, \shift_reg_1[7]_net_1\, 
        \shift_reg_1[8]_net_1\, \shift_reg_1[9]_net_1\, 
        \shift_reg_1[10]_net_1\, \shift_reg_1[11]_net_1\, 
        \shift_reg_1[12]_net_1\, \shift_reg_1[13]_net_1\, 
        \shift_reg_1[14]_net_1\, \shift_reg_0[0]_net_1\, 
        \shift_reg_0[1]_net_1\, \shift_reg_0[2]_net_1\, 
        \shift_reg_0[3]_net_1\, \shift_reg_0[4]_net_1\, 
        \shift_reg_0[5]_net_1\, \shift_reg_0[6]_net_1\, 
        \shift_reg_0[7]_net_1\, \shift_reg_0[8]_net_1\, 
        \shift_reg_0[9]_net_1\, \shift_reg_0[10]_net_1\, 
        \shift_reg_0[11]_net_1\, \shift_reg_0[12]_net_1\, 
        \shift_reg_0[13]_net_1\, \shift_reg_0[14]_net_1\, 
        \shift_reg_7[0]_net_1\, \shift_reg_7[1]_net_1\, 
        \shift_reg_7[2]_net_1\, \shift_reg_7[3]_net_1\, 
        \shift_reg_7[4]_net_1\, \shift_reg_7[5]_net_1\, 
        \shift_reg_7[6]_net_1\, \shift_reg_7[7]_net_1\, 
        \shift_reg_7[8]_net_1\, \shift_reg_7[9]_net_1\, 
        \shift_reg_7[10]_net_1\, \shift_reg_7[11]_net_1\, 
        \shift_reg_7[12]_net_1\, \shift_reg_7[13]_net_1\, 
        \shift_reg_7[14]_net_1\, \cnv_c\, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

    for all : SYNC_FF_1
	Use entity work.SYNC_FF_1(DEF_ARCH);
    for all : SYNC_FF
	Use entity work.SYNC_FF(DEF_ARCH);
begin 

    cnv_c <= \cnv_c\;

    \sample_bit_counter[2]\ : DFN1E0C0
      port map(D => N_13, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_6, Q => \sample_bit_counter[2]_net_1\);
    
    \shift_reg_0[1]\ : DFN1E1C0
      port map(D => \shift_reg_0[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[1]_net_1\);
    
    \cnv_cycle_counter_RNO_0[2]\ : AX1E
      port map(A => \cnv_cycle_counter[0]_net_1\, B => 
        \cnv_cycle_counter[1]_net_1\, C => 
        \cnv_cycle_counter[2]_net_1\, Y => 
        cnv_cycle_counter_n2_tz_i);
    
    \shift_reg_7[14]\ : DFN1E1C0
      port map(D => \shift_reg_7[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[14]_net_1\);
    
    \sample_6[13]\ : DFN1E1
      port map(D => \shift_reg_6[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(13));
    
    \sample_7[11]\ : DFN1E1
      port map(D => \shift_reg_7[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(11));
    
    \sample_0[3]\ : DFN1E1
      port map(D => \shift_reg_0[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(3));
    
    \shift_reg_6[12]\ : DFN1E1C0
      port map(D => \shift_reg_6[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[12]_net_1\);
    
    \sample_1[0]\ : DFN1E1
      port map(D => sdo_c(1), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(0));
    
    \sample_0[12]\ : DFN1E1
      port map(D => \shift_reg_0[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(12));
    
    \shift_reg_6[9]\ : DFN1E1C0
      port map(D => \shift_reg_6[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_6[9]_net_1\);
    
    \shift_reg_2[0]\ : DFN1E1C0
      port map(D => sdo_c(2), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_1[0]_net_1\, Q => 
        \shift_reg_2[0]_net_1\);
    
    \shift_reg_5[11]\ : DFN1E1C0
      port map(D => \shift_reg_5[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_5[11]_net_1\);
    
    cnv_s : DFN1C0
      port map(D => \cnv_s_RNO\, CLK => cnv_clk_c, CLR => 
        cnv_rstn_c, Q => \cnv_c\);
    
    \sample_6[11]\ : DFN1E1
      port map(D => \shift_reg_6[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(11));
    
    \sample_3[9]\ : DFN1E1
      port map(D => \shift_reg_3[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(9));
    
    \shift_reg_0[10]\ : DFN1E1C0
      port map(D => \shift_reg_0[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[10]_net_1\);
    
    \shift_reg_7[6]\ : DFN1E1C0
      port map(D => \shift_reg_7[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[6]_net_1\);
    
    \shift_reg_7[2]\ : DFN1E1C0
      port map(D => \shift_reg_7[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[2]_net_1\);
    
    \sample_2[6]\ : DFN1E1
      port map(D => \shift_reg_2[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(6));
    
    \cnv_cycle_counter[4]\ : DFN1C0
      port map(D => cnv_cycle_counter_n4, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[4]_net_1\);
    
    \cnv_cycle_counter_RNO[2]\ : NOR2
      port map(A => cnv_s_0_sqmuxa, B => 
        cnv_cycle_counter_n2_tz_i, Y => cnv_cycle_counter_n2);
    
    \sample_6[2]\ : DFN1E1
      port map(D => \shift_reg_6[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(2));
    
    \sample_7[5]\ : DFN1E1
      port map(D => \shift_reg_7[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(5));
    
    \shift_reg_5[6]\ : DFN1E1C0
      port map(D => \shift_reg_5[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[6]_net_1\);
    
    \shift_reg_0[14]\ : DFN1E1C0
      port map(D => \shift_reg_0[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[14]_net_1\);
    
    \shift_reg_1[7]\ : DFN1E1C0
      port map(D => \shift_reg_1[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[7]_net_1\);
    
    \sample_0[15]\ : DFN1E1
      port map(D => \shift_reg_0[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(15));
    
    \sample_2[4]\ : DFN1E1
      port map(D => \shift_reg_2[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(4));
    
    \sample_bit_counter_RNO[3]\ : XA1B
      port map(A => N_21, B => \sample_bit_counter[3]_net_1\, C
         => N_36, Y => N_15);
    
    \sample_1[6]\ : DFN1E1
      port map(D => \shift_reg_1[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(6));
    
    \cnv_cycle_counter_RNO[8]\ : XA1C
      port map(A => \cnv_cycle_counter[8]_net_1\, B => 
        cnv_cycle_counter_33_0, C => cnv_s_0_sqmuxa, Y => 
        cnv_cycle_counter_n8);
    
    \sample_2[14]\ : DFN1E1
      port map(D => \shift_reg_2[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(14));
    
    \sample_5[10]\ : DFN1E1
      port map(D => \shift_reg_5[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(10));
    
    \sample_2[0]\ : DFN1E1
      port map(D => sdo_c(2), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(0));
    
    \sample_5[1]\ : DFN1E1
      port map(D => \shift_reg_5[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(1));
    
    \shift_reg_4[13]\ : DFN1E1C0
      port map(D => \shift_reg_4[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[13]_net_1\);
    
    \cnv_cycle_counter_RNO[1]\ : XA1B
      port map(A => \cnv_cycle_counter[1]_net_1\, B => 
        \cnv_cycle_counter[0]_net_1\, C => cnv_s_0_sqmuxa, Y => 
        cnv_cycle_counter_n1);
    
    \shift_reg_7[5]\ : DFN1E1C0
      port map(D => \shift_reg_7[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[5]_net_1\);
    
    \sample_0[7]\ : DFN1E1
      port map(D => \shift_reg_0[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(7));
    
    \sample_0[13]\ : DFN1E1
      port map(D => \shift_reg_0[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(13));
    
    \shift_reg_1[10]\ : DFN1E1C0
      port map(D => \shift_reg_1[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_1[10]_net_1\);
    
    \sample_6[3]\ : DFN1E1
      port map(D => \shift_reg_6[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(3));
    
    \shift_reg_1[5]\ : DFN1E1C0
      port map(D => \shift_reg_1[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[5]_net_1\);
    
    \shift_reg_5[1]\ : DFN1E1C0
      port map(D => \shift_reg_5[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[1]_net_1\);
    
    \shift_reg_1[14]\ : DFN1E1C0
      port map(D => \shift_reg_1[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[14]_net_1\);
    
    cnv_done_RNO : OR2
      port map(A => cnv_sync_r_i_0, B => cnv_sync, Y => 
        cnv_done_1);
    
    \shift_reg_6[2]\ : DFN1E1C0
      port map(D => \shift_reg_6[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[2]_net_1\);
    
    \shift_reg_3[5]\ : DFN1E1C0
      port map(D => \shift_reg_3[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[5]_net_1\);
    
    cnv_done_RNI4H78 : AOI1B
      port map(A => \sample_bit_counter_0[0]_net_1\, B => 
        cnv_done_i, C => cnv_run_sync, Y => sample_bit_counter_n0);
    
    \sample_7[6]\ : DFN1E1
      port map(D => \shift_reg_7[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(6));
    
    \sample_7[10]\ : DFN1E1
      port map(D => \shift_reg_7[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(10));
    
    \sample_6[6]\ : DFN1E1
      port map(D => \shift_reg_6[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(6));
    
    \sample_0[11]\ : DFN1E1
      port map(D => \shift_reg_0[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(11));
    
    \shift_reg_0[0]\ : DFN1E1C0
      port map(D => sdo_c(0), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_0[0]_net_1\, Q => 
        \shift_reg_0[0]_net_1\);
    
    \sample_0[0]\ : DFN1E1
      port map(D => sdo_c(0), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(0));
    
    \sample_5[4]\ : DFN1E1
      port map(D => \shift_reg_5[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(4));
    
    \sample_7[9]\ : DFN1E1
      port map(D => \shift_reg_7[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(9));
    
    \sample_4[9]\ : DFN1E1
      port map(D => \shift_reg_4[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(9));
    
    \cnv_cycle_counter[6]\ : DFN1C0
      port map(D => cnv_cycle_counter_n6, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[6]_net_1\);
    
    \shift_reg_2[12]\ : DFN1E1C0
      port map(D => \shift_reg_2[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[12]_net_1\);
    
    \sample_bit_counter_1[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter_1[0]_net_1\);
    
    \sample_5[9]\ : DFN1E1
      port map(D => \shift_reg_5[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(9));
    
    \shift_reg_7[0]\ : DFN1E1C0
      port map(D => sdo_c(7), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[0]_net_1\);
    
    SYNC_FF_run : SYNC_FF_1
      port map(cnv_run_c => cnv_run_c, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, cnv_run_sync => cnv_run_sync);
    
    \shift_reg_1[1]\ : DFN1E1C0
      port map(D => \shift_reg_1[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[1]_net_1\);
    
    \shift_reg_3[9]\ : DFN1E1C0
      port map(D => \shift_reg_3[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_3[9]_net_1\);
    
    \sample_5[7]\ : DFN1E1
      port map(D => \shift_reg_5[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(7));
    
    \sample_bit_counter[5]\ : DFN1E0C0
      port map(D => N_19, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_6, Q => \sample_bit_counter[5]_net_1\);
    
    \sample_6[10]\ : DFN1E1
      port map(D => \shift_reg_6[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(10));
    
    \sample_3[12]\ : DFN1E1
      port map(D => \shift_reg_3[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(12));
    
    \shift_reg_3[6]\ : DFN1E1C0
      port map(D => \shift_reg_3[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[6]_net_1\);
    
    \sample_5[0]\ : DFN1E1
      port map(D => sdo_c(5), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(0));
    
    \sample_4[7]\ : DFN1E1
      port map(D => \shift_reg_4[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(7));
    
    \shift_reg_0[5]\ : DFN1E1C0
      port map(D => \shift_reg_0[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[5]_net_1\);
    
    \sample_bit_counter[4]\ : DFN1E0C0
      port map(D => N_17, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_6, Q => \sample_bit_counter[4]_net_1\);
    
    \sample_4[12]\ : DFN1E1
      port map(D => \shift_reg_4[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(12));
    
    \sample_2[7]\ : DFN1E1
      port map(D => \shift_reg_2[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(7));
    
    \shift_reg_7[8]\ : DFN1E1C0
      port map(D => \shift_reg_7[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[8]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \sample_bit_counter_RNID104[3]\ : NOR2B
      port map(A => \sample_bit_counter[3]_net_1\, B => N_21, Y
         => N_22);
    
    \shift_reg_0[3]\ : DFN1E1C0
      port map(D => \shift_reg_0[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[3]_net_1\);
    
    \sample_bit_counter_RNILHR2[2]\ : NOR2B
      port map(A => \sample_bit_counter[2]_net_1\, B => N_20, Y
         => N_21);
    
    \sample_bit_counter_RNIOIIL[5]\ : AO1A
      port map(A => N_36, B => \sample_bit_counter[5]_net_1\, C
         => N_30, Y => N_6);
    
    \shift_reg_6[11]\ : DFN1E1C0
      port map(D => \shift_reg_6[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[11]_net_1\);
    
    \sample_3[15]\ : DFN1E1
      port map(D => \shift_reg_3[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(15));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \shift_reg_3[8]\ : DFN1E1C0
      port map(D => \shift_reg_3[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[8]_net_1\);
    
    \shift_reg_4[10]\ : DFN1E1C0
      port map(D => \shift_reg_4[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[10]_net_1\);
    
    \sample_4[15]\ : DFN1E1
      port map(D => \shift_reg_4[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(15));
    
    \shift_reg_5[13]\ : DFN1E1C0
      port map(D => \shift_reg_5[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_5[13]_net_1\);
    
    \shift_reg_3[7]\ : DFN1E1C0
      port map(D => \shift_reg_3[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[7]_net_1\);
    
    \sample_0[2]\ : DFN1E1
      port map(D => \shift_reg_0[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(2));
    
    \cnv_cycle_counter_RNITOET[2]\ : OR2B
      port map(A => un2_cnv_run, B => cnv_run_c, Y => 
        cnv_s_0_sqmuxa);
    
    \shift_reg_4[14]\ : DFN1E1C0
      port map(D => \shift_reg_4[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[14]_net_1\);
    
    \sample_bit_counter_RNI8FD3[2]\ : NOR3
      port map(A => \sample_bit_counter[3]_net_1\, B => 
        \sample_bit_counter[2]_net_1\, C => 
        \sample_bit_counter[4]_net_1\, Y => 
        sample_bit_counterlde_i_a3_0_1);
    
    \sample_0[5]\ : DFN1E1
      port map(D => \shift_reg_0[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(5));
    
    \sample_3[13]\ : DFN1E1
      port map(D => \shift_reg_3[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(13));
    
    \sample_bit_counter_RNIVMI9_0[5]\ : CLKINT
      port map(A => \sample_bit_counter_RNIVMI9[5]_net_1\, Y => 
        sample_0_0_sqmuxa);
    
    \sample_2[5]\ : DFN1E1
      port map(D => \shift_reg_2[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(5));
    
    \shift_reg_2[5]\ : DFN1E1C0
      port map(D => \shift_reg_2[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[5]_net_1\);
    
    \sample_4[13]\ : DFN1E1
      port map(D => \shift_reg_4[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(13));
    
    \sample_3[1]\ : DFN1E1
      port map(D => \shift_reg_3[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(1));
    
    \sample_0[1]\ : DFN1E1
      port map(D => \shift_reg_0[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(1));
    
    \sample_0[10]\ : DFN1E1
      port map(D => \shift_reg_0[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(10));
    
    \shift_reg_0[2]\ : DFN1E1C0
      port map(D => \shift_reg_0[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[2]_net_1\);
    
    \sample_2[12]\ : DFN1E1
      port map(D => \shift_reg_2[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(12));
    
    \sample_6[0]\ : DFN1E1
      port map(D => sdo_c(6), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(0));
    
    \shift_reg_3[12]\ : DFN1E1C0
      port map(D => \shift_reg_3[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[12]_net_1\);
    
    \sample_val\ : DFN1C0
      port map(D => \sample_bit_counter_RNI0D96[5]_net_1\, CLK
         => HCLK_c, CLR => HRESETn_c, Q => sample_val);
    
    \cnv_cycle_counter_RNO[3]\ : NOR2
      port map(A => cnv_s_0_sqmuxa, B => 
        cnv_cycle_counter_n3_tz_i, Y => cnv_cycle_counter_n3);
    
    \sample_3[11]\ : DFN1E1
      port map(D => \shift_reg_3[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(11));
    
    \sample_0[9]\ : DFN1E1
      port map(D => \shift_reg_0[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(9));
    
    \shift_reg_5[8]\ : DFN1E1C0
      port map(D => \shift_reg_5[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[8]_net_1\);
    
    \sample_bit_counter_RNO[4]\ : XA1B
      port map(A => N_22, B => \sample_bit_counter[4]_net_1\, C
         => N_36, Y => N_17);
    
    \cnv_cycle_counter[3]\ : DFN1C0
      port map(D => cnv_cycle_counter_n3, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \sample_4[11]\ : DFN1E1
      port map(D => \shift_reg_4[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(11));
    
    \shift_reg_7[12]\ : DFN1E1C0
      port map(D => \shift_reg_7[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[12]_net_1\);
    
    \sample_6[7]\ : DFN1E1
      port map(D => \shift_reg_6[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(7));
    
    \sample_2[9]\ : DFN1E1
      port map(D => \shift_reg_2[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(9));
    
    \cnv_cycle_counter_RNO_0[8]\ : OR2B
      port map(A => cnv_cycle_counter_c6, B => 
        \cnv_cycle_counter[7]_net_1\, Y => cnv_cycle_counter_33_0);
    
    \shift_reg_6[1]\ : DFN1E1C0
      port map(D => \shift_reg_6[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[1]_net_1\);
    
    \shift_reg_7[7]\ : DFN1E1C0
      port map(D => \shift_reg_7[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[7]_net_1\);
    
    \sample_2[15]\ : DFN1E1
      port map(D => \shift_reg_2[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(15));
    
    \sample_bit_counter_0[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter_0[0]_net_1\);
    
    \shift_reg_6[3]\ : DFN1E1C0
      port map(D => \shift_reg_6[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[3]_net_1\);
    
    \sample_6[4]\ : DFN1E1
      port map(D => \shift_reg_6[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(4));
    
    \sample_4[3]\ : DFN1E1
      port map(D => \shift_reg_4[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(3));
    
    \sample_1[9]\ : DFN1E1
      port map(D => \shift_reg_1[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(9));
    
    \cnv_cycle_counter_RNO_0[4]\ : AX1E
      port map(A => \cnv_cycle_counter[3]_net_1\, B => 
        cnv_cycle_counter_c2, C => \cnv_cycle_counter[4]_net_1\, 
        Y => cnv_cycle_counter_n4_tz_i);
    
    \shift_reg_5[5]\ : DFN1E1C0
      port map(D => \shift_reg_5[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[5]_net_1\);
    
    \cnv_cycle_counter[7]\ : DFN1C0
      port map(D => cnv_cycle_counter_n7, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[7]_net_1\);
    
    \sample_1[14]\ : DFN1E1
      port map(D => \shift_reg_1[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(14));
    
    \shift_reg_2[11]\ : DFN1E1C0
      port map(D => \shift_reg_2[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[11]_net_1\);
    
    \shift_reg_7[3]\ : DFN1E1C0
      port map(D => \shift_reg_7[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[3]_net_1\);
    
    \shift_reg_5[10]\ : DFN1E1C0
      port map(D => \shift_reg_5[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_5[10]_net_1\);
    
    \shift_reg_3[4]\ : DFN1E1C0
      port map(D => \shift_reg_3[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[4]_net_1\);
    
    \sample_2[13]\ : DFN1E1
      port map(D => \shift_reg_2[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(13));
    
    \sample_bit_counter_RNI0D96[5]\ : NOR2
      port map(A => \sample_bit_counter[5]_net_1\, B => N_23, Y
         => \sample_bit_counter_RNI0D96[5]_net_1\);
    
    \sample_3[0]\ : DFN1E1
      port map(D => sdo_c(3), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(0));
    
    \shift_reg_0[12]\ : DFN1E1C0
      port map(D => \shift_reg_0[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[12]_net_1\);
    
    \sample_4[2]\ : DFN1E1
      port map(D => \shift_reg_4[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(2));
    
    \sample_bit_counter[1]\ : DFN1E0C0
      port map(D => N_11, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_6, Q => \sample_bit_counter[1]_net_1\);
    
    \shift_reg_5[14]\ : DFN1E1C0
      port map(D => \shift_reg_5[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[14]_net_1\);
    
    \sample_7[0]\ : DFN1E1
      port map(D => sdo_c(7), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(0));
    
    \sample_bit_counter_RNI28PC[2]\ : NOR3B
      port map(A => sample_bit_counterlde_i_a3_0_1, B => N_38, C
         => N_36, Y => N_30);
    
    \sample_2[3]\ : DFN1E1
      port map(D => \shift_reg_2[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(3));
    
    \sample_3[7]\ : DFN1E1
      port map(D => \shift_reg_3[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(7));
    
    \sample_7[1]\ : DFN1E1
      port map(D => \shift_reg_7[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(1));
    
    \sample_2[11]\ : DFN1E1
      port map(D => \shift_reg_2[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(11));
    
    cnv_sync_r : DFN1P0
      port map(D => cnv_sync_i, CLK => HCLK_c, PRE => HRESETn_c, 
        Q => cnv_sync_r_i_0);
    
    \cnv_cycle_counter_RNI6D3R[6]\ : NOR2A
      port map(A => \cnv_cycle_counter[6]_net_1\, B => 
        cnv_cycle_counter_c5, Y => cnv_cycle_counter_c6);
    
    \shift_reg_1[9]\ : DFN1E1C0
      port map(D => \shift_reg_1[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[9]_net_1\);
    
    \shift_reg_6[13]\ : DFN1E1C0
      port map(D => \shift_reg_6[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[13]_net_1\);
    
    \sample_6[1]\ : DFN1E1
      port map(D => \shift_reg_6[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(1));
    
    \shift_reg_0[8]\ : DFN1E1C0
      port map(D => \shift_reg_0[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[8]_net_1\);
    
    \sample_3[10]\ : DFN1E1
      port map(D => \shift_reg_3[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(10));
    
    \shift_reg_4[0]\ : DFN1E1C0
      port map(D => sdo_c(4), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_3[0]_net_1\, Q => 
        \shift_reg_4[0]_net_1\);
    
    SYNC_FF_cnv : SYNC_FF
      port map(cnv_c => \cnv_c\, HRESETn_c => HRESETn_c, HCLK_c
         => HCLK_c, cnv_sync => cnv_sync, cnv_sync_i => 
        cnv_sync_i);
    
    \shift_reg_2[2]\ : DFN1E1C0
      port map(D => \shift_reg_2[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[2]_net_1\);
    
    \sample_bit_counter_RNIU5N1_0[1]\ : NOR2
      port map(A => \sample_bit_counter[1]_net_1\, B => 
        \sample_bit_counter_0[0]_net_1\, Y => N_38);
    
    \shift_reg_1[3]\ : DFN1E1C0
      port map(D => \shift_reg_1[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[3]_net_1\);
    
    \shift_reg_1[12]\ : DFN1E1C0
      port map(D => \shift_reg_1[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[12]_net_1\);
    
    \sample_7[2]\ : DFN1E1
      port map(D => \shift_reg_7[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(2));
    
    \sample_4[10]\ : DFN1E1
      port map(D => \shift_reg_4[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(10));
    
    \sample_bit_counter_RNIU5N1[1]\ : NOR2B
      port map(A => \sample_bit_counter[1]_net_1\, B => 
        \sample_bit_counter_0[0]_net_1\, Y => N_20);
    
    \sample_3[8]\ : DFN1E1
      port map(D => \shift_reg_3[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(8));
    
    \shift_reg_3[3]\ : DFN1E1C0
      port map(D => \shift_reg_3[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[3]_net_1\);
    
    \shift_reg_1[8]\ : DFN1E1C0
      port map(D => \shift_reg_1[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[8]_net_1\);
    
    \sample_bit_counter_3[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter_3[0]_net_1\);
    
    \cnv_cycle_counter[8]\ : DFN1C0
      port map(D => cnv_cycle_counter_n8, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[8]_net_1\);
    
    \sample_bit_counter[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter[0]_net_1\);
    
    \sample_1[1]\ : DFN1E1
      port map(D => \shift_reg_1[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(1));
    
    \shift_reg_4[1]\ : DFN1E1C0
      port map(D => \shift_reg_4[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[1]_net_1\);
    
    \cnv_cycle_counter_RNO[0]\ : NOR2
      port map(A => \cnv_cycle_counter[0]_net_1\, B => 
        cnv_s_0_sqmuxa, Y => cnv_cycle_counter_n0);
    
    \sample_5[14]\ : DFN1E1
      port map(D => \shift_reg_5[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(14));
    
    \cnv_cycle_counter_RNIQQN7[8]\ : NOR2B
      port map(A => \cnv_cycle_counter[8]_net_1\, B => 
        \cnv_cycle_counter[4]_net_1\, Y => un2_cnv_runlto8_0);
    
    \shift_reg_3[1]\ : DFN1E1C0
      port map(D => \shift_reg_3[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[1]_net_1\);
    
    \shift_reg_2[8]\ : DFN1E1C0
      port map(D => \shift_reg_2[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[8]_net_1\);
    
    \sample_2[8]\ : DFN1E1
      port map(D => \shift_reg_2[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(8));
    
    \shift_reg_3[11]\ : DFN1E1C0
      port map(D => \shift_reg_3[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[11]_net_1\);
    
    \shift_reg_0[4]\ : DFN1E1C0
      port map(D => \shift_reg_0[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[4]_net_1\);
    
    \sample_4[5]\ : DFN1E1
      port map(D => \shift_reg_4[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(5));
    
    \sample_0[4]\ : DFN1E1
      port map(D => \shift_reg_0[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(4));
    
    \shift_reg_7[11]\ : DFN1E1C0
      port map(D => \shift_reg_7[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[11]_net_1\);
    
    \shift_reg_3[0]\ : DFN1E1C0
      port map(D => sdo_c(3), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_2[0]_net_1\, Q => 
        \shift_reg_3[0]_net_1\);
    
    \sample_3[4]\ : DFN1E1
      port map(D => \shift_reg_3[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(4));
    
    \sample_5[5]\ : DFN1E1
      port map(D => \shift_reg_5[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(5));
    
    \shift_reg_1[0]\ : DFN1E1C0
      port map(D => sdo_c(1), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_0[0]_net_1\, Q => 
        \shift_reg_1[0]_net_1\);
    
    \shift_reg_4[9]\ : DFN1E1C0
      port map(D => \shift_reg_4[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[9]_net_1\);
    
    \shift_reg_1[6]\ : DFN1E1C0
      port map(D => \shift_reg_1[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[6]_net_1\);
    
    \sample_4[1]\ : DFN1E1
      port map(D => \shift_reg_4[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(1));
    
    \shift_reg_2[9]\ : DFN1E1C0
      port map(D => \shift_reg_2[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[9]_net_1\);
    
    cnv_done_RNISIK7 : OR2B
      port map(A => cnv_run_sync, B => cnv_done_i, Y => N_36);
    
    \shift_reg_4[2]\ : DFN1E1C0
      port map(D => \shift_reg_4[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[2]_net_1\);
    
    \sample_7[8]\ : DFN1E1
      port map(D => \shift_reg_7[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(8));
    
    \sample_7[14]\ : DFN1E1
      port map(D => \shift_reg_7[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(14));
    
    \sample_2[10]\ : DFN1E1
      port map(D => \shift_reg_2[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(10));
    
    \shift_reg_6[10]\ : DFN1E1C0
      port map(D => \shift_reg_6[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[10]_net_1\);
    
    \shift_reg_3[2]\ : DFN1E1C0
      port map(D => \shift_reg_3[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[2]_net_1\);
    
    \shift_reg_4[12]\ : DFN1E1C0
      port map(D => \shift_reg_4[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[12]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \shift_reg_7[4]\ : DFN1E1C0
      port map(D => \shift_reg_7[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[4]_net_1\);
    
    \shift_reg_2[13]\ : DFN1E1C0
      port map(D => \shift_reg_2[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[13]_net_1\);
    
    \sample_6[5]\ : DFN1E1
      port map(D => \shift_reg_6[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(5));
    
    \shift_reg_6[14]\ : DFN1E1C0
      port map(D => \shift_reg_6[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[14]_net_1\);
    
    \cnv_cycle_counter_RNO[6]\ : XA1C
      port map(A => \cnv_cycle_counter[6]_net_1\, B => 
        cnv_cycle_counter_c5, C => cnv_s_0_sqmuxa, Y => 
        cnv_cycle_counter_n6);
    
    \sample_bit_counter_2[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter_2[0]_net_1\);
    
    \sample_5[2]\ : DFN1E1
      port map(D => \shift_reg_5[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(2));
    
    \sample_5[8]\ : DFN1E1
      port map(D => \shift_reg_5[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(8));
    
    \sample_1[12]\ : DFN1E1
      port map(D => \shift_reg_1[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(12));
    
    \shift_reg_2[6]\ : DFN1E1C0
      port map(D => \shift_reg_2[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[6]_net_1\);
    
    \shift_reg_0[11]\ : DFN1E1C0
      port map(D => \shift_reg_0[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[11]_net_1\);
    
    \sample_6[14]\ : DFN1E1
      port map(D => \shift_reg_6[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(14));
    
    cnv_s_RNO_0 : OA1C
      port map(A => \cnv_cycle_counter[6]_net_1\, B => 
        un3_cnv_runlt6, C => un3_cnv_runlto8_0, Y => un3_cnv_run);
    
    \shift_reg_4[8]\ : DFN1E1C0
      port map(D => \shift_reg_4[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[8]_net_1\);
    
    cnv_s_RNO_1 : AOI1
      port map(A => cnv_cycle_counter_c2, B => 
        \cnv_cycle_counter[3]_net_1\, C => un3_cnv_runlto5_0, Y
         => un3_cnv_runlt6);
    
    \cnv_cycle_counter[2]\ : DFN1C0
      port map(D => cnv_cycle_counter_n2, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[2]_net_1\);
    
    \sample_7[7]\ : DFN1E1
      port map(D => \shift_reg_7[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(7));
    
    \sample_3[5]\ : DFN1E1
      port map(D => \shift_reg_3[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(5));
    
    \shift_reg_7[1]\ : DFN1E1C0
      port map(D => \shift_reg_7[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[1]_net_1\);
    
    \sample_7[3]\ : DFN1E1
      port map(D => \shift_reg_7[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(3));
    
    \sample_3[6]\ : DFN1E1
      port map(D => \shift_reg_3[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(6));
    
    \cnv_cycle_counter_RNO[5]\ : XA1B
      port map(A => \cnv_cycle_counter[5]_net_1\, B => 
        cnv_cycle_counter_c4, C => cnv_s_0_sqmuxa, Y => 
        cnv_cycle_counter_n5);
    
    \shift_reg_5[9]\ : DFN1E1C0
      port map(D => \shift_reg_5[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[9]_net_1\);
    
    \shift_reg_4[6]\ : DFN1E1C0
      port map(D => \shift_reg_4[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[6]_net_1\);
    
    \shift_reg_1[4]\ : DFN1E1C0
      port map(D => \shift_reg_1[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[4]_net_1\);
    
    \cnv_cycle_counter_RNIPQN7[5]\ : NOR2B
      port map(A => \cnv_cycle_counter[5]_net_1\, B => 
        \cnv_cycle_counter[6]_net_1\, Y => un2_cnv_runlto8_1);
    
    \shift_reg_4[5]\ : DFN1E1C0
      port map(D => \shift_reg_4[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[5]_net_1\);
    
    \sample_2[1]\ : DFN1E1
      port map(D => \shift_reg_2[0]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(1));
    
    \sample_1[15]\ : DFN1E1
      port map(D => \shift_reg_1[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(15));
    
    sck : DFN1P0
      port map(D => \sample_bit_counter_i[0]\, CLK => HCLK_c, PRE
         => HRESETn_c, Q => sck_c);
    
    \shift_reg_6[8]\ : DFN1E1C0
      port map(D => \shift_reg_6[7]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_6[8]_net_1\);
    
    \shift_reg_5[4]\ : DFN1E1C0
      port map(D => \shift_reg_5[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[4]_net_1\);
    
    \cnv_cycle_counter_RNO[4]\ : NOR2
      port map(A => cnv_s_0_sqmuxa, B => 
        cnv_cycle_counter_n4_tz_i, Y => cnv_cycle_counter_n4);
    
    \sample_bit_counter_RNO[2]\ : XA1B
      port map(A => N_20, B => \sample_bit_counter[2]_net_1\, C
         => N_36, Y => N_13);
    
    \sample_5[6]\ : DFN1E1
      port map(D => \shift_reg_5[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(6));
    
    \sample_bit_counter_4[0]\ : DFN1E0C0
      port map(D => sample_bit_counter_n0, CLK => HCLK_c, CLR => 
        HRESETn_c, E => N_6, Q => \sample_bit_counter_4[0]_net_1\);
    
    \shift_reg_0[6]\ : DFN1E1C0
      port map(D => \shift_reg_0[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[6]_net_1\);
    
    \sample_1[3]\ : DFN1E1
      port map(D => \shift_reg_1[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(3));
    
    \cnv_cycle_counter_RNIONJB[1]\ : NOR3C
      port map(A => \cnv_cycle_counter[0]_net_1\, B => 
        \cnv_cycle_counter[1]_net_1\, C => 
        \cnv_cycle_counter[2]_net_1\, Y => cnv_cycle_counter_c2);
    
    \shift_reg_5[3]\ : DFN1E1C0
      port map(D => \shift_reg_5[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[3]_net_1\);
    
    \sample_3[2]\ : DFN1E1
      port map(D => \shift_reg_3[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(2));
    
    \sample_5[3]\ : DFN1E1
      port map(D => \shift_reg_5[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(3));
    
    \shift_reg_1[11]\ : DFN1E1C0
      port map(D => \shift_reg_1[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[11]_net_1\);
    
    \sample_bit_counter_RNO[5]\ : NOR2
      port map(A => N_36, B => N_23, Y => N_19);
    
    \cnv_cycle_counter[5]\ : DFN1C0
      port map(D => cnv_cycle_counter_n5, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[5]_net_1\);
    
    \sample_1[7]\ : DFN1E1
      port map(D => \shift_reg_1[6]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(7));
    
    \sample_1[13]\ : DFN1E1
      port map(D => \shift_reg_1[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(13));
    
    sck_RNO : INV
      port map(A => \sample_bit_counter_0[0]_net_1\, Y => 
        \sample_bit_counter_i[0]\);
    
    \shift_reg_5[2]\ : DFN1E1C0
      port map(D => \shift_reg_5[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[2]_net_1\);
    
    \sample_bit_counter_RNO[1]\ : NOR3
      port map(A => N_38, B => N_36, C => N_20, Y => N_11);
    
    \sample_6[8]\ : DFN1E1
      port map(D => \shift_reg_6[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(8));
    
    \sample_1[2]\ : DFN1E1
      port map(D => \shift_reg_1[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(2));
    
    \sample_bit_counter_RNI6L45[4]\ : OR2B
      port map(A => \sample_bit_counter[4]_net_1\, B => N_22, Y
         => N_23);
    
    \cnv_cycle_counter_RNIKD3R[2]\ : OR3C
      port map(A => un2_cnv_runlto8_1, B => un2_cnv_runlto8_0, C
         => un2_cnv_runlto8_2, Y => un2_cnv_run);
    
    \sample_0[8]\ : DFN1E1
      port map(D => \shift_reg_0[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(8));
    
    \sample_0[14]\ : DFN1E1
      port map(D => \shift_reg_0[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(14));
    
    \sample_5[12]\ : DFN1E1
      port map(D => \shift_reg_5[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(12));
    
    \shift_reg_0[9]\ : DFN1E1C0
      port map(D => \shift_reg_0[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[9]_net_1\);
    
    \sample_bit_counter_RNIVMI9[5]\ : NOR2B
      port map(A => \sample_bit_counter_RNI0D96[5]_net_1\, B => 
        HRESETn_c, Y => \sample_bit_counter_RNIVMI9[5]_net_1\);
    
    \sample_1[11]\ : DFN1E1
      port map(D => \shift_reg_1[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(11));
    
    \shift_reg_5[7]\ : DFN1E1C0
      port map(D => \shift_reg_5[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_5[7]_net_1\);
    
    \sample_0[6]\ : DFN1E1
      port map(D => \shift_reg_0[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_0(6));
    
    \shift_reg_2[10]\ : DFN1E1C0
      port map(D => \shift_reg_2[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[10]_net_1\);
    
    \shift_reg_5[12]\ : DFN1E1C0
      port map(D => \shift_reg_5[11]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_5[12]_net_1\);
    
    \shift_reg_3[13]\ : DFN1E1C0
      port map(D => \shift_reg_3[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[13]_net_1\);
    
    cnv_done : DFN1P0
      port map(D => cnv_done_1, CLK => HCLK_c, PRE => HRESETn_c, 
        Q => cnv_done_i);
    
    \shift_reg_2[1]\ : DFN1E1C0
      port map(D => \shift_reg_2[0]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[1]_net_1\);
    
    \sample_7[4]\ : DFN1E1
      port map(D => \shift_reg_7[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(4));
    
    \sample_4[6]\ : DFN1E1
      port map(D => \shift_reg_4[5]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(6));
    
    \shift_reg_1[2]\ : DFN1E1C0
      port map(D => \shift_reg_1[1]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[2]_net_1\);
    
    cnv_s_RNO_3 : OR2
      port map(A => \cnv_cycle_counter[4]_net_1\, B => 
        \cnv_cycle_counter[5]_net_1\, Y => un3_cnv_runlto5_0);
    
    \shift_reg_7[13]\ : DFN1E1C0
      port map(D => \shift_reg_7[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[13]_net_1\);
    
    \shift_reg_2[14]\ : DFN1E1C0
      port map(D => \shift_reg_2[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_2[14]_net_1\);
    
    \cnv_cycle_counter_RNIDIBJ[4]\ : NOR3C
      port map(A => \cnv_cycle_counter[3]_net_1\, B => 
        cnv_cycle_counter_c2, C => \cnv_cycle_counter[4]_net_1\, 
        Y => cnv_cycle_counter_c4);
    
    \shift_reg_6[5]\ : DFN1E1C0
      port map(D => \shift_reg_6[4]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[5]_net_1\);
    
    \sample_4[8]\ : DFN1E1
      port map(D => \shift_reg_4[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(8));
    
    \sample_5[15]\ : DFN1E1
      port map(D => \shift_reg_5[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(15));
    
    \shift_reg_2[3]\ : DFN1E1C0
      port map(D => \shift_reg_2[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[3]_net_1\);
    
    cnv_s_RNO : OA1A
      port map(A => un2_cnv_run, B => un3_cnv_run, C => cnv_run_c, 
        Y => \cnv_s_RNO\);
    
    \shift_reg_6[0]\ : DFN1E1C0
      port map(D => sdo_c(6), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_4[0]_net_1\, Q => 
        \shift_reg_6[0]_net_1\);
    
    \cnv_cycle_counter[0]\ : DFN1C0
      port map(D => cnv_cycle_counter_n0, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[0]_net_1\);
    
    \shift_reg_2[7]\ : DFN1E1C0
      port map(D => \shift_reg_2[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[7]_net_1\);
    
    \shift_reg_6[4]\ : DFN1E1C0
      port map(D => \shift_reg_6[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_4[0]_net_1\, Q
         => \shift_reg_6[4]_net_1\);
    
    \shift_reg_2[4]\ : DFN1E1C0
      port map(D => \shift_reg_2[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_2[4]_net_1\);
    
    \sample_6[9]\ : DFN1E1
      port map(D => \shift_reg_6[8]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(9));
    
    \shift_reg_4[4]\ : DFN1E1C0
      port map(D => \shift_reg_4[3]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[4]_net_1\);
    
    \sample_7[12]\ : DFN1E1
      port map(D => \shift_reg_7[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(12));
    
    \cnv_cycle_counter_RNIPF7N[5]\ : OR2B
      port map(A => cnv_cycle_counter_c4, B => 
        \cnv_cycle_counter[5]_net_1\, Y => cnv_cycle_counter_c5);
    
    \shift_reg_4[3]\ : DFN1E1C0
      port map(D => \shift_reg_4[2]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[3]_net_1\);
    
    \shift_reg_4[11]\ : DFN1E1C0
      port map(D => \shift_reg_4[10]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[11]_net_1\);
    
    \sample_bit_counter[3]\ : DFN1E0C0
      port map(D => N_15, CLK => HCLK_c, CLR => HRESETn_c, E => 
        N_6, Q => \sample_bit_counter[3]_net_1\);
    
    \cnv_cycle_counter_RNI1OJB[2]\ : OA1
      port map(A => \cnv_cycle_counter[2]_net_1\, B => 
        \cnv_cycle_counter[3]_net_1\, C => 
        \cnv_cycle_counter[7]_net_1\, Y => un2_cnv_runlto8_2);
    
    \sample_5[13]\ : DFN1E1
      port map(D => \shift_reg_5[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(13));
    
    \shift_reg_0[7]\ : DFN1E1C0
      port map(D => \shift_reg_0[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[7]_net_1\);
    
    cnv_s_RNO_2 : OR2
      port map(A => \cnv_cycle_counter[8]_net_1\, B => 
        \cnv_cycle_counter[7]_net_1\, Y => un3_cnv_runlto8_0);
    
    \shift_reg_0[13]\ : DFN1E1C0
      port map(D => \shift_reg_0[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_0[0]_net_1\, Q
         => \shift_reg_0[13]_net_1\);
    
    \sample_2[2]\ : DFN1E1
      port map(D => \shift_reg_2[1]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_2(2));
    
    \sample_1[8]\ : DFN1E1
      port map(D => \shift_reg_1[7]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(8));
    
    \sample_1[5]\ : DFN1E1
      port map(D => \shift_reg_1[4]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(5));
    
    \sample_6[12]\ : DFN1E1
      port map(D => \shift_reg_6[11]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(12));
    
    \cnv_cycle_counter_RNO[7]\ : XA1B
      port map(A => \cnv_cycle_counter[7]_net_1\, B => 
        cnv_cycle_counter_c6, C => cnv_s_0_sqmuxa, Y => 
        cnv_cycle_counter_n7);
    
    \sample_7[15]\ : DFN1E1
      port map(D => \shift_reg_7[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(15));
    
    \sample_4[0]\ : DFN1E1
      port map(D => sdo_c(4), CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(0));
    
    \shift_reg_5[0]\ : DFN1E1C0
      port map(D => sdo_c(5), CLK => HCLK_c, CLR => HRESETn_c, E
         => \sample_bit_counter_3[0]_net_1\, Q => 
        \shift_reg_5[0]_net_1\);
    
    \sample_3[3]\ : DFN1E1
      port map(D => \shift_reg_3[2]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(3));
    
    \sample_5[11]\ : DFN1E1
      port map(D => \shift_reg_5[10]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_5(11));
    
    \shift_reg_4[7]\ : DFN1E1C0
      port map(D => \shift_reg_4[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_3[0]_net_1\, Q
         => \shift_reg_4[7]_net_1\);
    
    \shift_reg_6[6]\ : DFN1E1C0
      port map(D => \shift_reg_6[5]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_6[6]_net_1\);
    
    \sample_4[4]\ : DFN1E1
      port map(D => \shift_reg_4[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(4));
    
    \sample_6[15]\ : DFN1E1
      port map(D => \shift_reg_6[14]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_6(15));
    
    \shift_reg_3[10]\ : DFN1E1C0
      port map(D => \shift_reg_3[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[10]_net_1\);
    
    \sample_1[10]\ : DFN1E1
      port map(D => \shift_reg_1[9]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(10));
    
    \sample_3[14]\ : DFN1E1
      port map(D => \shift_reg_3[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_3(14));
    
    \sample_7[13]\ : DFN1E1
      port map(D => \shift_reg_7[12]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_7(13));
    
    \shift_reg_7[9]\ : DFN1E1C0
      port map(D => \shift_reg_7[8]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[9]_net_1\);
    
    \sample_1[4]\ : DFN1E1
      port map(D => \shift_reg_1[3]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_1(4));
    
    \cnv_cycle_counter_RNO_0[3]\ : XNOR2
      port map(A => cnv_cycle_counter_c2, B => 
        \cnv_cycle_counter[3]_net_1\, Y => 
        cnv_cycle_counter_n3_tz_i);
    
    \cnv_cycle_counter[1]\ : DFN1C0
      port map(D => cnv_cycle_counter_n1, CLK => cnv_clk_c, CLR
         => cnv_rstn_c, Q => \cnv_cycle_counter[1]_net_1\);
    
    \shift_reg_7[10]\ : DFN1E1C0
      port map(D => \shift_reg_7[9]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_7[10]_net_1\);
    
    \sample_4[14]\ : DFN1E1
      port map(D => \shift_reg_4[13]_net_1\, CLK => HCLK_c, E => 
        sample_0_0_sqmuxa, Q => sample_4(14));
    
    \shift_reg_6[7]\ : DFN1E1C0
      port map(D => \shift_reg_6[6]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter[0]_net_1\, Q => 
        \shift_reg_6[7]_net_1\);
    
    \shift_reg_3[14]\ : DFN1E1C0
      port map(D => \shift_reg_3[13]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_2[0]_net_1\, Q
         => \shift_reg_3[14]_net_1\);
    
    \shift_reg_1[13]\ : DFN1E1C0
      port map(D => \shift_reg_1[12]_net_1\, CLK => HCLK_c, CLR
         => HRESETn_c, E => \sample_bit_counter_1[0]_net_1\, Q
         => \shift_reg_1[13]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_top_lfr_wf_picker_ip is

    port( nb_snapshot_param            : in    std_logic_vector(10 downto 0);
          delta_f2_f0                  : in    std_logic_vector(9 downto 0);
          delta_snapshot               : in    std_logic_vector(15 downto 0);
          delta_f2_f1                  : in    std_logic_vector(9 downto 0);
          status_new_err               : out   std_logic_vector(3 downto 0);
          hwdata_c                     : out   std_logic_vector(31 downto 0);
          addr_data_f0                 : in    std_logic_vector(31 downto 0);
          addr_data_f1                 : in    std_logic_vector(31 downto 0);
          addr_data_f2                 : in    std_logic_vector(31 downto 0);
          addr_data_f3                 : in    std_logic_vector(31 downto 0);
          status_full                  : out   std_logic_vector(3 downto 0);
          status_full_err              : out   std_logic_vector(3 downto 0);
          nb_burst_available           : in    std_logic_vector(10 downto 0);
          haddr_c                      : out   std_logic_vector(31 downto 0);
          AHB_Master_In_c_3            : in    std_logic;
          AHB_Master_In_c_0            : in    std_logic;
          AHB_Master_In_c_4            : in    std_logic;
          AHB_Master_In_c_5            : in    std_logic;
          hsize_c                      : out   std_logic_vector(1 downto 0);
          htrans_c                     : out   std_logic_vector(1 downto 0);
          hburst_c                     : out   std_logic_vector(2 downto 0);
          status_full_ack              : in    std_logic_vector(3 downto 0);
          sdo_c                        : in    std_logic_vector(7 downto 0);
          coarse_time_0_c              : in    std_logic;
          enable_f0                    : in    std_logic;
          data_shaping_R0              : in    std_logic;
          data_shaping_R0_0            : in    std_logic;
          burst_f0                     : in    std_logic;
          data_shaping_R1              : in    std_logic;
          data_shaping_R1_0            : in    std_logic;
          enable_f1                    : in    std_logic;
          burst_f1                     : in    std_logic;
          enable_f2                    : in    std_logic;
          burst_f2                     : in    std_logic;
          enable_f3                    : in    std_logic;
          N_43                         : out   std_logic;
          IdlePhase_RNI03G71           : out   std_logic;
          hwrite_c                     : out   std_logic;
          lpp_top_lfr_wf_picker_ip_GND : in    std_logic;
          lpp_top_lfr_wf_picker_ip_VCC : in    std_logic;
          cnv_run_c                    : in    std_logic;
          sck_c                        : out   std_logic;
          cnv_c                        : out   std_logic;
          cnv_clk_c                    : in    std_logic;
          cnv_rstn_c                   : in    std_logic;
          data_shaping_SP0             : in    std_logic;
          data_shaping_SP1             : in    std_logic;
          HRESETn_c                    : in    std_logic;
          HCLK_c                       : in    std_logic
        );

end lpp_top_lfr_wf_picker_ip;

architecture DEF_ARCH of lpp_top_lfr_wf_picker_ip is 

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IIR_CEL_CTRLR_v2
    port( sample_filter_v2_out_0   : out   std_logic;
          sample_filter_v2_out_1   : out   std_logic;
          sample_filter_v2_out_2   : out   std_logic;
          sample_filter_v2_out_3   : out   std_logic;
          sample_filter_v2_out_4   : out   std_logic;
          sample_filter_v2_out_5   : out   std_logic;
          sample_filter_v2_out_6   : out   std_logic;
          sample_filter_v2_out_7   : out   std_logic;
          sample_filter_v2_out_8   : out   std_logic;
          sample_filter_v2_out_9   : out   std_logic;
          sample_filter_v2_out_10  : out   std_logic;
          sample_filter_v2_out_11  : out   std_logic;
          sample_filter_v2_out_12  : out   std_logic;
          sample_filter_v2_out_13  : out   std_logic;
          sample_filter_v2_out_14  : out   std_logic;
          sample_filter_v2_out_15  : out   std_logic;
          sample_filter_v2_out_18  : out   std_logic;
          sample_filter_v2_out_19  : out   std_logic;
          sample_filter_v2_out_20  : out   std_logic;
          sample_filter_v2_out_21  : out   std_logic;
          sample_filter_v2_out_22  : out   std_logic;
          sample_filter_v2_out_23  : out   std_logic;
          sample_filter_v2_out_24  : out   std_logic;
          sample_filter_v2_out_25  : out   std_logic;
          sample_filter_v2_out_26  : out   std_logic;
          sample_filter_v2_out_27  : out   std_logic;
          sample_filter_v2_out_28  : out   std_logic;
          sample_filter_v2_out_29  : out   std_logic;
          sample_filter_v2_out_30  : out   std_logic;
          sample_filter_v2_out_31  : out   std_logic;
          sample_filter_v2_out_32  : out   std_logic;
          sample_filter_v2_out_33  : out   std_logic;
          sample_filter_v2_out_36  : out   std_logic;
          sample_filter_v2_out_37  : out   std_logic;
          sample_filter_v2_out_38  : out   std_logic;
          sample_filter_v2_out_39  : out   std_logic;
          sample_filter_v2_out_40  : out   std_logic;
          sample_filter_v2_out_41  : out   std_logic;
          sample_filter_v2_out_42  : out   std_logic;
          sample_filter_v2_out_43  : out   std_logic;
          sample_filter_v2_out_44  : out   std_logic;
          sample_filter_v2_out_45  : out   std_logic;
          sample_filter_v2_out_46  : out   std_logic;
          sample_filter_v2_out_47  : out   std_logic;
          sample_filter_v2_out_48  : out   std_logic;
          sample_filter_v2_out_49  : out   std_logic;
          sample_filter_v2_out_50  : out   std_logic;
          sample_filter_v2_out_51  : out   std_logic;
          sample_filter_v2_out_54  : out   std_logic;
          sample_filter_v2_out_55  : out   std_logic;
          sample_filter_v2_out_56  : out   std_logic;
          sample_filter_v2_out_57  : out   std_logic;
          sample_filter_v2_out_58  : out   std_logic;
          sample_filter_v2_out_59  : out   std_logic;
          sample_filter_v2_out_60  : out   std_logic;
          sample_filter_v2_out_61  : out   std_logic;
          sample_filter_v2_out_62  : out   std_logic;
          sample_filter_v2_out_63  : out   std_logic;
          sample_filter_v2_out_64  : out   std_logic;
          sample_filter_v2_out_65  : out   std_logic;
          sample_filter_v2_out_66  : out   std_logic;
          sample_filter_v2_out_67  : out   std_logic;
          sample_filter_v2_out_68  : out   std_logic;
          sample_filter_v2_out_69  : out   std_logic;
          sample_filter_v2_out_90  : out   std_logic;
          sample_filter_v2_out_91  : out   std_logic;
          sample_filter_v2_out_92  : out   std_logic;
          sample_filter_v2_out_93  : out   std_logic;
          sample_filter_v2_out_94  : out   std_logic;
          sample_filter_v2_out_95  : out   std_logic;
          sample_filter_v2_out_96  : out   std_logic;
          sample_filter_v2_out_97  : out   std_logic;
          sample_filter_v2_out_98  : out   std_logic;
          sample_filter_v2_out_99  : out   std_logic;
          sample_filter_v2_out_100 : out   std_logic;
          sample_filter_v2_out_101 : out   std_logic;
          sample_filter_v2_out_102 : out   std_logic;
          sample_filter_v2_out_103 : out   std_logic;
          sample_filter_v2_out_104 : out   std_logic;
          sample_filter_v2_out_105 : out   std_logic;
          sample_filter_v2_out_108 : out   std_logic;
          sample_filter_v2_out_126 : out   std_logic;
          sample_filter_v2_out_109 : out   std_logic;
          sample_filter_v2_out_127 : out   std_logic;
          sample_filter_v2_out_110 : out   std_logic;
          sample_filter_v2_out_128 : out   std_logic;
          sample_filter_v2_out_111 : out   std_logic;
          sample_filter_v2_out_129 : out   std_logic;
          sample_filter_v2_out_112 : out   std_logic;
          sample_filter_v2_out_130 : out   std_logic;
          sample_filter_v2_out_113 : out   std_logic;
          sample_filter_v2_out_131 : out   std_logic;
          sample_filter_v2_out_114 : out   std_logic;
          sample_filter_v2_out_132 : out   std_logic;
          sample_filter_v2_out_115 : out   std_logic;
          sample_filter_v2_out_133 : out   std_logic;
          sample_filter_v2_out_116 : out   std_logic;
          sample_filter_v2_out_134 : out   std_logic;
          sample_filter_v2_out_117 : out   std_logic;
          sample_filter_v2_out_135 : out   std_logic;
          sample_filter_v2_out_118 : out   std_logic;
          sample_filter_v2_out_136 : out   std_logic;
          sample_filter_v2_out_119 : out   std_logic;
          sample_filter_v2_out_137 : out   std_logic;
          sample_filter_v2_out_120 : out   std_logic;
          sample_filter_v2_out_138 : out   std_logic;
          sample_filter_v2_out_121 : out   std_logic;
          sample_filter_v2_out_139 : out   std_logic;
          sample_filter_v2_out_122 : out   std_logic;
          sample_filter_v2_out_140 : out   std_logic;
          sample_filter_v2_out_123 : out   std_logic;
          sample_filter_v2_out_141 : out   std_logic;
          sample_6                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_5                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_2                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_0                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_1                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_3                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_4                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          sample_7                 : in    std_logic_vector(15 downto 0) := (others => 'U');
          IIR_CEL_CTRLR_v2_VCC     : in    std_logic := 'U';
          IIR_CEL_CTRLR_v2_GND     : in    std_logic := 'U';
          HRESETn_c                : in    std_logic := 'U';
          HCLK_c                   : in    std_logic := 'U';
          sample_filter_v2_out_val : out   std_logic;
          sample_val_delay         : in    std_logic := 'U'
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component Downsampling_6_16_256
    port( sample_f1          : in    std_logic_vector(111 downto 80) := (others => 'U');
          sample_f1_wdata_95 : in    std_logic := 'U';
          sample_f1_wdata_94 : in    std_logic := 'U';
          sample_f1_wdata_93 : in    std_logic := 'U';
          sample_f1_wdata_92 : in    std_logic := 'U';
          sample_f1_wdata_91 : in    std_logic := 'U';
          sample_f1_wdata_90 : in    std_logic := 'U';
          sample_f1_wdata_89 : in    std_logic := 'U';
          sample_f1_wdata_88 : in    std_logic := 'U';
          sample_f1_wdata_87 : in    std_logic := 'U';
          sample_f1_wdata_86 : in    std_logic := 'U';
          sample_f1_wdata_85 : in    std_logic := 'U';
          sample_f1_wdata_84 : in    std_logic := 'U';
          sample_f1_wdata_83 : in    std_logic := 'U';
          sample_f1_wdata_82 : in    std_logic := 'U';
          sample_f1_wdata_81 : in    std_logic := 'U';
          sample_f1_wdata_80 : in    std_logic := 'U';
          sample_f1_wdata_79 : in    std_logic := 'U';
          sample_f1_wdata_78 : in    std_logic := 'U';
          sample_f1_wdata_77 : in    std_logic := 'U';
          sample_f1_wdata_76 : in    std_logic := 'U';
          sample_f1_wdata_75 : in    std_logic := 'U';
          sample_f1_wdata_74 : in    std_logic := 'U';
          sample_f1_wdata_73 : in    std_logic := 'U';
          sample_f1_wdata_72 : in    std_logic := 'U';
          sample_f1_wdata_71 : in    std_logic := 'U';
          sample_f1_wdata_70 : in    std_logic := 'U';
          sample_f1_wdata_69 : in    std_logic := 'U';
          sample_f1_wdata_68 : in    std_logic := 'U';
          sample_f1_wdata_67 : in    std_logic := 'U';
          sample_f1_wdata_66 : in    std_logic := 'U';
          sample_f1_wdata_65 : in    std_logic := 'U';
          sample_f1_wdata_64 : in    std_logic := 'U';
          sample_f1_wdata_63 : in    std_logic := 'U';
          sample_f1_wdata_62 : in    std_logic := 'U';
          sample_f1_wdata_61 : in    std_logic := 'U';
          sample_f1_wdata_60 : in    std_logic := 'U';
          sample_f1_wdata_59 : in    std_logic := 'U';
          sample_f1_wdata_58 : in    std_logic := 'U';
          sample_f1_wdata_57 : in    std_logic := 'U';
          sample_f1_wdata_56 : in    std_logic := 'U';
          sample_f1_wdata_55 : in    std_logic := 'U';
          sample_f1_wdata_54 : in    std_logic := 'U';
          sample_f1_wdata_53 : in    std_logic := 'U';
          sample_f1_wdata_52 : in    std_logic := 'U';
          sample_f1_wdata_51 : in    std_logic := 'U';
          sample_f1_wdata_50 : in    std_logic := 'U';
          sample_f1_wdata_49 : in    std_logic := 'U';
          sample_f1_wdata_48 : in    std_logic := 'U';
          sample_f1_wdata_15 : in    std_logic := 'U';
          sample_f1_wdata_14 : in    std_logic := 'U';
          sample_f1_wdata_13 : in    std_logic := 'U';
          sample_f1_wdata_12 : in    std_logic := 'U';
          sample_f1_wdata_11 : in    std_logic := 'U';
          sample_f1_wdata_10 : in    std_logic := 'U';
          sample_f1_wdata_9  : in    std_logic := 'U';
          sample_f1_wdata_8  : in    std_logic := 'U';
          sample_f1_wdata_7  : in    std_logic := 'U';
          sample_f1_wdata_6  : in    std_logic := 'U';
          sample_f1_wdata_5  : in    std_logic := 'U';
          sample_f1_wdata_4  : in    std_logic := 'U';
          sample_f1_wdata_3  : in    std_logic := 'U';
          sample_f1_wdata_2  : in    std_logic := 'U';
          sample_f1_wdata_1  : in    std_logic := 'U';
          sample_f1_wdata_0  : in    std_logic := 'U';
          sample_f3_wdata    : out   std_logic_vector(95 downto 0);
          sample_f1_val      : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          sample_f3_val      : out   std_logic;
          HRESETn_c          : in    std_logic := 'U';
          sample_f1_val_0    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Downsampling_6_16_96
    port( sample_f0             : in    std_logic_vector(111 downto 80) := (others => 'U');
          sample_f0_wdata_95    : in    std_logic := 'U';
          sample_f0_wdata_94    : in    std_logic := 'U';
          sample_f0_wdata_93    : in    std_logic := 'U';
          sample_f0_wdata_92    : in    std_logic := 'U';
          sample_f0_wdata_91    : in    std_logic := 'U';
          sample_f0_wdata_90    : in    std_logic := 'U';
          sample_f0_wdata_89    : in    std_logic := 'U';
          sample_f0_wdata_88    : in    std_logic := 'U';
          sample_f0_wdata_87    : in    std_logic := 'U';
          sample_f0_wdata_86    : in    std_logic := 'U';
          sample_f0_wdata_85    : in    std_logic := 'U';
          sample_f0_wdata_84    : in    std_logic := 'U';
          sample_f0_wdata_83    : in    std_logic := 'U';
          sample_f0_wdata_82    : in    std_logic := 'U';
          sample_f0_wdata_81    : in    std_logic := 'U';
          sample_f0_wdata_80    : in    std_logic := 'U';
          sample_f0_wdata_79    : in    std_logic := 'U';
          sample_f0_wdata_78    : in    std_logic := 'U';
          sample_f0_wdata_77    : in    std_logic := 'U';
          sample_f0_wdata_76    : in    std_logic := 'U';
          sample_f0_wdata_75    : in    std_logic := 'U';
          sample_f0_wdata_74    : in    std_logic := 'U';
          sample_f0_wdata_73    : in    std_logic := 'U';
          sample_f0_wdata_72    : in    std_logic := 'U';
          sample_f0_wdata_71    : in    std_logic := 'U';
          sample_f0_wdata_70    : in    std_logic := 'U';
          sample_f0_wdata_69    : in    std_logic := 'U';
          sample_f0_wdata_68    : in    std_logic := 'U';
          sample_f0_wdata_67    : in    std_logic := 'U';
          sample_f0_wdata_66    : in    std_logic := 'U';
          sample_f0_wdata_65    : in    std_logic := 'U';
          sample_f0_wdata_64    : in    std_logic := 'U';
          sample_f0_wdata_63    : in    std_logic := 'U';
          sample_f0_wdata_62    : in    std_logic := 'U';
          sample_f0_wdata_61    : in    std_logic := 'U';
          sample_f0_wdata_60    : in    std_logic := 'U';
          sample_f0_wdata_59    : in    std_logic := 'U';
          sample_f0_wdata_58    : in    std_logic := 'U';
          sample_f0_wdata_57    : in    std_logic := 'U';
          sample_f0_wdata_56    : in    std_logic := 'U';
          sample_f0_wdata_55    : in    std_logic := 'U';
          sample_f0_wdata_54    : in    std_logic := 'U';
          sample_f0_wdata_53    : in    std_logic := 'U';
          sample_f0_wdata_52    : in    std_logic := 'U';
          sample_f0_wdata_51    : in    std_logic := 'U';
          sample_f0_wdata_50    : in    std_logic := 'U';
          sample_f0_wdata_49    : in    std_logic := 'U';
          sample_f0_wdata_48    : in    std_logic := 'U';
          sample_f0_wdata_15    : in    std_logic := 'U';
          sample_f0_wdata_14    : in    std_logic := 'U';
          sample_f0_wdata_13    : in    std_logic := 'U';
          sample_f0_wdata_12    : in    std_logic := 'U';
          sample_f0_wdata_11    : in    std_logic := 'U';
          sample_f0_wdata_10    : in    std_logic := 'U';
          sample_f0_wdata_9     : in    std_logic := 'U';
          sample_f0_wdata_8     : in    std_logic := 'U';
          sample_f0_wdata_7     : in    std_logic := 'U';
          sample_f0_wdata_6     : in    std_logic := 'U';
          sample_f0_wdata_5     : in    std_logic := 'U';
          sample_f0_wdata_4     : in    std_logic := 'U';
          sample_f0_wdata_3     : in    std_logic := 'U';
          sample_f0_wdata_2     : in    std_logic := 'U';
          sample_f0_wdata_1     : in    std_logic := 'U';
          sample_f0_wdata_0     : in    std_logic := 'U';
          sample_f2_wdata       : out   std_logic_vector(95 downto 0);
          sample_f0_val         : in    std_logic := 'U';
          sample_f0_val_1       : in    std_logic := 'U';
          HRESETn_c             : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U';
          sample_f2_val         : out   std_logic;
          sample_f0_val_0       : in    std_logic := 'U';
          sample_out_0_sqmuxa_1 : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component lpp_waveform
    port( status_full_ack    : in    std_logic_vector(3 downto 0) := (others => 'U');
          hburst_c           : out   std_logic_vector(2 downto 0);
          htrans_c           : out   std_logic_vector(1 downto 0);
          hsize_c            : out   std_logic_vector(1 downto 0);
          AHB_Master_In_c_5  : in    std_logic := 'U';
          AHB_Master_In_c_4  : in    std_logic := 'U';
          AHB_Master_In_c_0  : in    std_logic := 'U';
          AHB_Master_In_c_3  : in    std_logic := 'U';
          haddr_c            : out   std_logic_vector(31 downto 0);
          nb_burst_available : in    std_logic_vector(10 downto 0) := (others => 'U');
          status_full_err    : out   std_logic_vector(3 downto 0);
          status_full        : out   std_logic_vector(3 downto 0);
          addr_data_f3       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f2       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f1       : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f0       : in    std_logic_vector(31 downto 0) := (others => 'U');
          hwdata_c           : out   std_logic_vector(31 downto 0);
          status_new_err     : out   std_logic_vector(3 downto 0);
          sample_f3_wdata    : in    std_logic_vector(95 downto 0) := (others => 'U');
          sample_f2_wdata    : in    std_logic_vector(95 downto 0) := (others => 'U');
          sample_f1_15       : in    std_logic := 'U';
          sample_f1_47       : in    std_logic := 'U';
          sample_f1_14       : in    std_logic := 'U';
          sample_f1_46       : in    std_logic := 'U';
          sample_f1_13       : in    std_logic := 'U';
          sample_f1_45       : in    std_logic := 'U';
          sample_f1_12       : in    std_logic := 'U';
          sample_f1_44       : in    std_logic := 'U';
          sample_f1_60       : in    std_logic := 'U';
          sample_f1_59       : in    std_logic := 'U';
          sample_f1_58       : in    std_logic := 'U';
          sample_f1_57       : in    std_logic := 'U';
          sample_f1_56       : in    std_logic := 'U';
          sample_f1_55       : in    std_logic := 'U';
          sample_f1_54       : in    std_logic := 'U';
          sample_f1_53       : in    std_logic := 'U';
          sample_f1_52       : in    std_logic := 'U';
          sample_f1_51       : in    std_logic := 'U';
          sample_f1_50       : in    std_logic := 'U';
          sample_f1_49       : in    std_logic := 'U';
          sample_f1_48       : in    std_logic := 'U';
          sample_f1_4        : in    std_logic := 'U';
          sample_f1_36       : in    std_logic := 'U';
          sample_f1_3        : in    std_logic := 'U';
          sample_f1_35       : in    std_logic := 'U';
          sample_f1_2        : in    std_logic := 'U';
          sample_f1_34       : in    std_logic := 'U';
          sample_f1_1        : in    std_logic := 'U';
          sample_f1_33       : in    std_logic := 'U';
          sample_f1_0        : in    std_logic := 'U';
          sample_f1_32       : in    std_logic := 'U';
          sample_f1_63       : in    std_logic := 'U';
          sample_f1_62       : in    std_logic := 'U';
          sample_f1_61       : in    std_logic := 'U';
          sample_f1_11       : in    std_logic := 'U';
          sample_f1_43       : in    std_logic := 'U';
          sample_f1_10       : in    std_logic := 'U';
          sample_f1_42       : in    std_logic := 'U';
          sample_f1_9        : in    std_logic := 'U';
          sample_f1_41       : in    std_logic := 'U';
          sample_f1_8        : in    std_logic := 'U';
          sample_f1_40       : in    std_logic := 'U';
          sample_f1_7        : in    std_logic := 'U';
          sample_f1_39       : in    std_logic := 'U';
          sample_f1_6        : in    std_logic := 'U';
          sample_f1_38       : in    std_logic := 'U';
          sample_f1_5        : in    std_logic := 'U';
          sample_f1_37       : in    std_logic := 'U';
          sample_f1_wdata_0  : in    std_logic := 'U';
          sample_f1_wdata_1  : in    std_logic := 'U';
          sample_f1_wdata_2  : in    std_logic := 'U';
          sample_f1_wdata_3  : in    std_logic := 'U';
          sample_f1_wdata_4  : in    std_logic := 'U';
          sample_f1_wdata_5  : in    std_logic := 'U';
          sample_f1_wdata_6  : in    std_logic := 'U';
          sample_f1_wdata_7  : in    std_logic := 'U';
          sample_f1_wdata_8  : in    std_logic := 'U';
          sample_f1_wdata_9  : in    std_logic := 'U';
          sample_f1_wdata_10 : in    std_logic := 'U';
          sample_f1_wdata_11 : in    std_logic := 'U';
          sample_f1_wdata_12 : in    std_logic := 'U';
          sample_f1_wdata_13 : in    std_logic := 'U';
          sample_f1_wdata_14 : in    std_logic := 'U';
          sample_f1_wdata_15 : in    std_logic := 'U';
          sample_f1_wdata_48 : in    std_logic := 'U';
          sample_f1_wdata_49 : in    std_logic := 'U';
          sample_f1_wdata_50 : in    std_logic := 'U';
          sample_f1_wdata_51 : in    std_logic := 'U';
          sample_f1_wdata_52 : in    std_logic := 'U';
          sample_f1_wdata_53 : in    std_logic := 'U';
          sample_f1_wdata_54 : in    std_logic := 'U';
          sample_f1_wdata_55 : in    std_logic := 'U';
          sample_f1_wdata_56 : in    std_logic := 'U';
          sample_f1_wdata_57 : in    std_logic := 'U';
          sample_f1_wdata_58 : in    std_logic := 'U';
          sample_f1_wdata_59 : in    std_logic := 'U';
          sample_f1_wdata_60 : in    std_logic := 'U';
          sample_f1_wdata_61 : in    std_logic := 'U';
          sample_f1_wdata_62 : in    std_logic := 'U';
          sample_f1_wdata_63 : in    std_logic := 'U';
          sample_f1_wdata_64 : in    std_logic := 'U';
          sample_f1_wdata_65 : in    std_logic := 'U';
          sample_f1_wdata_66 : in    std_logic := 'U';
          sample_f1_wdata_67 : in    std_logic := 'U';
          sample_f1_wdata_68 : in    std_logic := 'U';
          sample_f1_wdata_69 : in    std_logic := 'U';
          sample_f1_wdata_70 : in    std_logic := 'U';
          sample_f1_wdata_71 : in    std_logic := 'U';
          sample_f1_wdata_72 : in    std_logic := 'U';
          sample_f1_wdata_73 : in    std_logic := 'U';
          sample_f1_wdata_74 : in    std_logic := 'U';
          sample_f1_wdata_75 : in    std_logic := 'U';
          sample_f1_wdata_76 : in    std_logic := 'U';
          sample_f1_wdata_77 : in    std_logic := 'U';
          sample_f1_wdata_78 : in    std_logic := 'U';
          sample_f1_wdata_79 : in    std_logic := 'U';
          sample_f1_wdata_80 : in    std_logic := 'U';
          sample_f1_wdata_81 : in    std_logic := 'U';
          sample_f1_wdata_82 : in    std_logic := 'U';
          sample_f1_wdata_83 : in    std_logic := 'U';
          sample_f1_wdata_84 : in    std_logic := 'U';
          sample_f1_wdata_85 : in    std_logic := 'U';
          sample_f1_wdata_86 : in    std_logic := 'U';
          sample_f1_wdata_87 : in    std_logic := 'U';
          sample_f1_wdata_88 : in    std_logic := 'U';
          sample_f1_wdata_89 : in    std_logic := 'U';
          sample_f1_wdata_90 : in    std_logic := 'U';
          sample_f1_wdata_91 : in    std_logic := 'U';
          sample_f1_wdata_92 : in    std_logic := 'U';
          sample_f1_wdata_93 : in    std_logic := 'U';
          sample_f1_wdata_94 : in    std_logic := 'U';
          sample_f1_wdata_95 : in    std_logic := 'U';
          sample_f0_15       : in    std_logic := 'U';
          sample_f0_47       : in    std_logic := 'U';
          sample_f0_14       : in    std_logic := 'U';
          sample_f0_46       : in    std_logic := 'U';
          sample_f0_13       : in    std_logic := 'U';
          sample_f0_45       : in    std_logic := 'U';
          sample_f0_12       : in    std_logic := 'U';
          sample_f0_44       : in    std_logic := 'U';
          sample_f0_60       : in    std_logic := 'U';
          sample_f0_59       : in    std_logic := 'U';
          sample_f0_58       : in    std_logic := 'U';
          sample_f0_57       : in    std_logic := 'U';
          sample_f0_56       : in    std_logic := 'U';
          sample_f0_55       : in    std_logic := 'U';
          sample_f0_54       : in    std_logic := 'U';
          sample_f0_53       : in    std_logic := 'U';
          sample_f0_52       : in    std_logic := 'U';
          sample_f0_51       : in    std_logic := 'U';
          sample_f0_50       : in    std_logic := 'U';
          sample_f0_49       : in    std_logic := 'U';
          sample_f0_48       : in    std_logic := 'U';
          sample_f0_4        : in    std_logic := 'U';
          sample_f0_36       : in    std_logic := 'U';
          sample_f0_3        : in    std_logic := 'U';
          sample_f0_35       : in    std_logic := 'U';
          sample_f0_2        : in    std_logic := 'U';
          sample_f0_34       : in    std_logic := 'U';
          sample_f0_1        : in    std_logic := 'U';
          sample_f0_33       : in    std_logic := 'U';
          sample_f0_0        : in    std_logic := 'U';
          sample_f0_32       : in    std_logic := 'U';
          sample_f0_63       : in    std_logic := 'U';
          sample_f0_62       : in    std_logic := 'U';
          sample_f0_61       : in    std_logic := 'U';
          sample_f0_11       : in    std_logic := 'U';
          sample_f0_43       : in    std_logic := 'U';
          sample_f0_10       : in    std_logic := 'U';
          sample_f0_42       : in    std_logic := 'U';
          sample_f0_9        : in    std_logic := 'U';
          sample_f0_41       : in    std_logic := 'U';
          sample_f0_8        : in    std_logic := 'U';
          sample_f0_40       : in    std_logic := 'U';
          sample_f0_7        : in    std_logic := 'U';
          sample_f0_39       : in    std_logic := 'U';
          sample_f0_6        : in    std_logic := 'U';
          sample_f0_38       : in    std_logic := 'U';
          sample_f0_5        : in    std_logic := 'U';
          sample_f0_37       : in    std_logic := 'U';
          sample_f0_wdata_0  : in    std_logic := 'U';
          sample_f0_wdata_1  : in    std_logic := 'U';
          sample_f0_wdata_2  : in    std_logic := 'U';
          sample_f0_wdata_3  : in    std_logic := 'U';
          sample_f0_wdata_4  : in    std_logic := 'U';
          sample_f0_wdata_5  : in    std_logic := 'U';
          sample_f0_wdata_6  : in    std_logic := 'U';
          sample_f0_wdata_7  : in    std_logic := 'U';
          sample_f0_wdata_8  : in    std_logic := 'U';
          sample_f0_wdata_9  : in    std_logic := 'U';
          sample_f0_wdata_10 : in    std_logic := 'U';
          sample_f0_wdata_11 : in    std_logic := 'U';
          sample_f0_wdata_12 : in    std_logic := 'U';
          sample_f0_wdata_13 : in    std_logic := 'U';
          sample_f0_wdata_14 : in    std_logic := 'U';
          sample_f0_wdata_15 : in    std_logic := 'U';
          sample_f0_wdata_48 : in    std_logic := 'U';
          sample_f0_wdata_49 : in    std_logic := 'U';
          sample_f0_wdata_50 : in    std_logic := 'U';
          sample_f0_wdata_51 : in    std_logic := 'U';
          sample_f0_wdata_52 : in    std_logic := 'U';
          sample_f0_wdata_53 : in    std_logic := 'U';
          sample_f0_wdata_54 : in    std_logic := 'U';
          sample_f0_wdata_55 : in    std_logic := 'U';
          sample_f0_wdata_56 : in    std_logic := 'U';
          sample_f0_wdata_57 : in    std_logic := 'U';
          sample_f0_wdata_58 : in    std_logic := 'U';
          sample_f0_wdata_59 : in    std_logic := 'U';
          sample_f0_wdata_60 : in    std_logic := 'U';
          sample_f0_wdata_61 : in    std_logic := 'U';
          sample_f0_wdata_62 : in    std_logic := 'U';
          sample_f0_wdata_63 : in    std_logic := 'U';
          sample_f0_wdata_64 : in    std_logic := 'U';
          sample_f0_wdata_65 : in    std_logic := 'U';
          sample_f0_wdata_66 : in    std_logic := 'U';
          sample_f0_wdata_67 : in    std_logic := 'U';
          sample_f0_wdata_68 : in    std_logic := 'U';
          sample_f0_wdata_69 : in    std_logic := 'U';
          sample_f0_wdata_70 : in    std_logic := 'U';
          sample_f0_wdata_71 : in    std_logic := 'U';
          sample_f0_wdata_72 : in    std_logic := 'U';
          sample_f0_wdata_73 : in    std_logic := 'U';
          sample_f0_wdata_74 : in    std_logic := 'U';
          sample_f0_wdata_75 : in    std_logic := 'U';
          sample_f0_wdata_76 : in    std_logic := 'U';
          sample_f0_wdata_77 : in    std_logic := 'U';
          sample_f0_wdata_78 : in    std_logic := 'U';
          sample_f0_wdata_79 : in    std_logic := 'U';
          sample_f0_wdata_80 : in    std_logic := 'U';
          sample_f0_wdata_81 : in    std_logic := 'U';
          sample_f0_wdata_82 : in    std_logic := 'U';
          sample_f0_wdata_83 : in    std_logic := 'U';
          sample_f0_wdata_84 : in    std_logic := 'U';
          sample_f0_wdata_85 : in    std_logic := 'U';
          sample_f0_wdata_86 : in    std_logic := 'U';
          sample_f0_wdata_87 : in    std_logic := 'U';
          sample_f0_wdata_88 : in    std_logic := 'U';
          sample_f0_wdata_89 : in    std_logic := 'U';
          sample_f0_wdata_90 : in    std_logic := 'U';
          sample_f0_wdata_91 : in    std_logic := 'U';
          sample_f0_wdata_92 : in    std_logic := 'U';
          sample_f0_wdata_93 : in    std_logic := 'U';
          sample_f0_wdata_94 : in    std_logic := 'U';
          sample_f0_wdata_95 : in    std_logic := 'U';
          delta_f2_f1        : in    std_logic_vector(9 downto 0) := (others => 'U');
          delta_snapshot     : in    std_logic_vector(15 downto 0) := (others => 'U');
          delta_f2_f0        : in    std_logic_vector(9 downto 0) := (others => 'U');
          nb_snapshot_param  : in    std_logic_vector(10 downto 0) := (others => 'U');
          hwrite_c           : out   std_logic;
          IdlePhase_RNI03G71 : out   std_logic;
          N_43               : out   std_logic;
          lpp_waveform_GND   : in    std_logic := 'U';
          lpp_waveform_VCC   : in    std_logic := 'U';
          sample_f3_val      : in    std_logic := 'U';
          enable_f3          : in    std_logic := 'U';
          burst_f2           : in    std_logic := 'U';
          enable_f2          : in    std_logic := 'U';
          sample_f1_val_0    : in    std_logic := 'U';
          burst_f1           : in    std_logic := 'U';
          enable_f1          : in    std_logic := 'U';
          data_shaping_R1_0  : in    std_logic := 'U';
          data_shaping_R1    : in    std_logic := 'U';
          burst_f0           : in    std_logic := 'U';
          data_shaping_R0_0  : in    std_logic := 'U';
          data_shaping_R0    : in    std_logic := 'U';
          enable_f0          : in    std_logic := 'U';
          coarse_time_0_c    : in    std_logic := 'U';
          sample_f2_val      : in    std_logic := 'U';
          sample_f0_val_0    : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          HRESETn_c          : in    std_logic := 'U'
        );
  end component;

  component Downsampling_8_16_4
    port( sample_f0_0                   : out   std_logic;
          sample_f0_1                   : out   std_logic;
          sample_f0_2                   : out   std_logic;
          sample_f0_3                   : out   std_logic;
          sample_f0_4                   : out   std_logic;
          sample_f0_5                   : out   std_logic;
          sample_f0_6                   : out   std_logic;
          sample_f0_7                   : out   std_logic;
          sample_f0_8                   : out   std_logic;
          sample_f0_9                   : out   std_logic;
          sample_f0_10                  : out   std_logic;
          sample_f0_11                  : out   std_logic;
          sample_f0_12                  : out   std_logic;
          sample_f0_13                  : out   std_logic;
          sample_f0_14                  : out   std_logic;
          sample_f0_15                  : out   std_logic;
          sample_f0_32                  : out   std_logic;
          sample_f0_33                  : out   std_logic;
          sample_f0_34                  : out   std_logic;
          sample_f0_35                  : out   std_logic;
          sample_f0_36                  : out   std_logic;
          sample_f0_37                  : out   std_logic;
          sample_f0_38                  : out   std_logic;
          sample_f0_39                  : out   std_logic;
          sample_f0_40                  : out   std_logic;
          sample_f0_41                  : out   std_logic;
          sample_f0_42                  : out   std_logic;
          sample_f0_43                  : out   std_logic;
          sample_f0_44                  : out   std_logic;
          sample_f0_45                  : out   std_logic;
          sample_f0_46                  : out   std_logic;
          sample_f0_47                  : out   std_logic;
          sample_f0_48                  : out   std_logic;
          sample_f0_49                  : out   std_logic;
          sample_f0_50                  : out   std_logic;
          sample_f0_51                  : out   std_logic;
          sample_f0_52                  : out   std_logic;
          sample_f0_53                  : out   std_logic;
          sample_f0_54                  : out   std_logic;
          sample_f0_55                  : out   std_logic;
          sample_f0_56                  : out   std_logic;
          sample_f0_57                  : out   std_logic;
          sample_f0_58                  : out   std_logic;
          sample_f0_59                  : out   std_logic;
          sample_f0_60                  : out   std_logic;
          sample_f0_61                  : out   std_logic;
          sample_f0_62                  : out   std_logic;
          sample_f0_63                  : out   std_logic;
          sample_data_shaping_out_0     : in    std_logic := 'U';
          sample_data_shaping_out_1     : in    std_logic := 'U';
          sample_data_shaping_out_2     : in    std_logic := 'U';
          sample_data_shaping_out_3     : in    std_logic := 'U';
          sample_data_shaping_out_4     : in    std_logic := 'U';
          sample_data_shaping_out_5     : in    std_logic := 'U';
          sample_data_shaping_out_6     : in    std_logic := 'U';
          sample_data_shaping_out_7     : in    std_logic := 'U';
          sample_data_shaping_out_8     : in    std_logic := 'U';
          sample_data_shaping_out_9     : in    std_logic := 'U';
          sample_data_shaping_out_10    : in    std_logic := 'U';
          sample_data_shaping_out_11    : in    std_logic := 'U';
          sample_data_shaping_out_12    : in    std_logic := 'U';
          sample_data_shaping_out_13    : in    std_logic := 'U';
          sample_data_shaping_out_14    : in    std_logic := 'U';
          sample_data_shaping_out_15    : in    std_logic := 'U';
          sample_data_shaping_out_18    : in    std_logic := 'U';
          sample_data_shaping_out_19    : in    std_logic := 'U';
          sample_data_shaping_out_20    : in    std_logic := 'U';
          sample_data_shaping_out_21    : in    std_logic := 'U';
          sample_data_shaping_out_22    : in    std_logic := 'U';
          sample_data_shaping_out_23    : in    std_logic := 'U';
          sample_data_shaping_out_24    : in    std_logic := 'U';
          sample_data_shaping_out_25    : in    std_logic := 'U';
          sample_data_shaping_out_26    : in    std_logic := 'U';
          sample_data_shaping_out_27    : in    std_logic := 'U';
          sample_data_shaping_out_28    : in    std_logic := 'U';
          sample_data_shaping_out_29    : in    std_logic := 'U';
          sample_data_shaping_out_30    : in    std_logic := 'U';
          sample_data_shaping_out_31    : in    std_logic := 'U';
          sample_data_shaping_out_32    : in    std_logic := 'U';
          sample_data_shaping_out_33    : in    std_logic := 'U';
          sample_data_shaping_out_36    : in    std_logic := 'U';
          sample_data_shaping_out_37    : in    std_logic := 'U';
          sample_data_shaping_out_38    : in    std_logic := 'U';
          sample_data_shaping_out_39    : in    std_logic := 'U';
          sample_data_shaping_out_40    : in    std_logic := 'U';
          sample_data_shaping_out_41    : in    std_logic := 'U';
          sample_data_shaping_out_42    : in    std_logic := 'U';
          sample_data_shaping_out_43    : in    std_logic := 'U';
          sample_data_shaping_out_44    : in    std_logic := 'U';
          sample_data_shaping_out_45    : in    std_logic := 'U';
          sample_data_shaping_out_46    : in    std_logic := 'U';
          sample_data_shaping_out_47    : in    std_logic := 'U';
          sample_data_shaping_out_48    : in    std_logic := 'U';
          sample_data_shaping_out_49    : in    std_logic := 'U';
          sample_data_shaping_out_50    : in    std_logic := 'U';
          sample_data_shaping_out_51    : in    std_logic := 'U';
          sample_data_shaping_out_54    : in    std_logic := 'U';
          sample_data_shaping_out_55    : in    std_logic := 'U';
          sample_data_shaping_out_56    : in    std_logic := 'U';
          sample_data_shaping_out_57    : in    std_logic := 'U';
          sample_data_shaping_out_58    : in    std_logic := 'U';
          sample_data_shaping_out_59    : in    std_logic := 'U';
          sample_data_shaping_out_60    : in    std_logic := 'U';
          sample_data_shaping_out_61    : in    std_logic := 'U';
          sample_data_shaping_out_62    : in    std_logic := 'U';
          sample_data_shaping_out_63    : in    std_logic := 'U';
          sample_data_shaping_out_64    : in    std_logic := 'U';
          sample_data_shaping_out_65    : in    std_logic := 'U';
          sample_data_shaping_out_66    : in    std_logic := 'U';
          sample_data_shaping_out_67    : in    std_logic := 'U';
          sample_data_shaping_out_68    : in    std_logic := 'U';
          sample_data_shaping_out_69    : in    std_logic := 'U';
          sample_data_shaping_out_90    : in    std_logic := 'U';
          sample_data_shaping_out_91    : in    std_logic := 'U';
          sample_data_shaping_out_92    : in    std_logic := 'U';
          sample_data_shaping_out_93    : in    std_logic := 'U';
          sample_data_shaping_out_94    : in    std_logic := 'U';
          sample_data_shaping_out_95    : in    std_logic := 'U';
          sample_data_shaping_out_96    : in    std_logic := 'U';
          sample_data_shaping_out_97    : in    std_logic := 'U';
          sample_data_shaping_out_98    : in    std_logic := 'U';
          sample_data_shaping_out_99    : in    std_logic := 'U';
          sample_data_shaping_out_100   : in    std_logic := 'U';
          sample_data_shaping_out_101   : in    std_logic := 'U';
          sample_data_shaping_out_102   : in    std_logic := 'U';
          sample_data_shaping_out_103   : in    std_logic := 'U';
          sample_data_shaping_out_104   : in    std_logic := 'U';
          sample_data_shaping_out_105   : in    std_logic := 'U';
          sample_data_shaping_out_108   : in    std_logic := 'U';
          sample_data_shaping_out_109   : in    std_logic := 'U';
          sample_data_shaping_out_110   : in    std_logic := 'U';
          sample_data_shaping_out_111   : in    std_logic := 'U';
          sample_data_shaping_out_112   : in    std_logic := 'U';
          sample_data_shaping_out_113   : in    std_logic := 'U';
          sample_data_shaping_out_114   : in    std_logic := 'U';
          sample_data_shaping_out_115   : in    std_logic := 'U';
          sample_data_shaping_out_116   : in    std_logic := 'U';
          sample_data_shaping_out_117   : in    std_logic := 'U';
          sample_data_shaping_out_118   : in    std_logic := 'U';
          sample_data_shaping_out_119   : in    std_logic := 'U';
          sample_data_shaping_out_120   : in    std_logic := 'U';
          sample_data_shaping_out_121   : in    std_logic := 'U';
          sample_data_shaping_out_122   : in    std_logic := 'U';
          sample_data_shaping_out_123   : in    std_logic := 'U';
          sample_data_shaping_out_126   : in    std_logic := 'U';
          sample_data_shaping_out_127   : in    std_logic := 'U';
          sample_data_shaping_out_128   : in    std_logic := 'U';
          sample_data_shaping_out_129   : in    std_logic := 'U';
          sample_data_shaping_out_130   : in    std_logic := 'U';
          sample_data_shaping_out_131   : in    std_logic := 'U';
          sample_data_shaping_out_132   : in    std_logic := 'U';
          sample_data_shaping_out_133   : in    std_logic := 'U';
          sample_data_shaping_out_134   : in    std_logic := 'U';
          sample_data_shaping_out_135   : in    std_logic := 'U';
          sample_data_shaping_out_136   : in    std_logic := 'U';
          sample_data_shaping_out_137   : in    std_logic := 'U';
          sample_data_shaping_out_138   : in    std_logic := 'U';
          sample_data_shaping_out_139   : in    std_logic := 'U';
          sample_data_shaping_out_140   : in    std_logic := 'U';
          sample_data_shaping_out_141   : in    std_logic := 'U';
          sample_f0_wdata_95            : out   std_logic;
          sample_f0_wdata_94            : out   std_logic;
          sample_f0_wdata_93            : out   std_logic;
          sample_f0_wdata_92            : out   std_logic;
          sample_f0_wdata_91            : out   std_logic;
          sample_f0_wdata_90            : out   std_logic;
          sample_f0_wdata_89            : out   std_logic;
          sample_f0_wdata_88            : out   std_logic;
          sample_f0_wdata_87            : out   std_logic;
          sample_f0_wdata_86            : out   std_logic;
          sample_f0_wdata_85            : out   std_logic;
          sample_f0_wdata_84            : out   std_logic;
          sample_f0_wdata_83            : out   std_logic;
          sample_f0_wdata_82            : out   std_logic;
          sample_f0_wdata_81            : out   std_logic;
          sample_f0_wdata_80            : out   std_logic;
          sample_f0_wdata_79            : out   std_logic;
          sample_f0_wdata_78            : out   std_logic;
          sample_f0_wdata_77            : out   std_logic;
          sample_f0_wdata_76            : out   std_logic;
          sample_f0_wdata_75            : out   std_logic;
          sample_f0_wdata_74            : out   std_logic;
          sample_f0_wdata_73            : out   std_logic;
          sample_f0_wdata_72            : out   std_logic;
          sample_f0_wdata_71            : out   std_logic;
          sample_f0_wdata_70            : out   std_logic;
          sample_f0_wdata_69            : out   std_logic;
          sample_f0_wdata_68            : out   std_logic;
          sample_f0_wdata_67            : out   std_logic;
          sample_f0_wdata_66            : out   std_logic;
          sample_f0_wdata_65            : out   std_logic;
          sample_f0_wdata_64            : out   std_logic;
          sample_f0_wdata_63            : out   std_logic;
          sample_f0_wdata_62            : out   std_logic;
          sample_f0_wdata_61            : out   std_logic;
          sample_f0_wdata_60            : out   std_logic;
          sample_f0_wdata_59            : out   std_logic;
          sample_f0_wdata_58            : out   std_logic;
          sample_f0_wdata_57            : out   std_logic;
          sample_f0_wdata_56            : out   std_logic;
          sample_f0_wdata_55            : out   std_logic;
          sample_f0_wdata_54            : out   std_logic;
          sample_f0_wdata_53            : out   std_logic;
          sample_f0_wdata_52            : out   std_logic;
          sample_f0_wdata_51            : out   std_logic;
          sample_f0_wdata_50            : out   std_logic;
          sample_f0_wdata_49            : out   std_logic;
          sample_f0_wdata_48            : out   std_logic;
          sample_f0_wdata_15            : out   std_logic;
          sample_f0_wdata_14            : out   std_logic;
          sample_f0_wdata_13            : out   std_logic;
          sample_f0_wdata_12            : out   std_logic;
          sample_f0_wdata_11            : out   std_logic;
          sample_f0_wdata_10            : out   std_logic;
          sample_f0_wdata_9             : out   std_logic;
          sample_f0_wdata_8             : out   std_logic;
          sample_f0_wdata_7             : out   std_logic;
          sample_f0_wdata_6             : out   std_logic;
          sample_f0_wdata_5             : out   std_logic;
          sample_f0_wdata_4             : out   std_logic;
          sample_f0_wdata_3             : out   std_logic;
          sample_f0_wdata_2             : out   std_logic;
          sample_f0_wdata_1             : out   std_logic;
          sample_f0_wdata_0             : out   std_logic;
          sample_data_shaping_out_val   : in    std_logic := 'U';
          sample_f0_val                 : out   std_logic;
          sample_data_shaping_out_val_0 : in    std_logic := 'U';
          sample_f0_val_0               : out   std_logic;
          HRESETn_c                     : in    std_logic := 'U';
          HCLK_c                        : in    std_logic := 'U';
          sample_f0_val_1               : out   std_logic
        );
  end component;

  component Downsampling_8_16_6
    port( sample_f0_0           : in    std_logic := 'U';
          sample_f0_1           : in    std_logic := 'U';
          sample_f0_2           : in    std_logic := 'U';
          sample_f0_3           : in    std_logic := 'U';
          sample_f0_4           : in    std_logic := 'U';
          sample_f0_5           : in    std_logic := 'U';
          sample_f0_6           : in    std_logic := 'U';
          sample_f0_7           : in    std_logic := 'U';
          sample_f0_8           : in    std_logic := 'U';
          sample_f0_9           : in    std_logic := 'U';
          sample_f0_10          : in    std_logic := 'U';
          sample_f0_11          : in    std_logic := 'U';
          sample_f0_12          : in    std_logic := 'U';
          sample_f0_13          : in    std_logic := 'U';
          sample_f0_14          : in    std_logic := 'U';
          sample_f0_15          : in    std_logic := 'U';
          sample_f0_32          : in    std_logic := 'U';
          sample_f0_33          : in    std_logic := 'U';
          sample_f0_34          : in    std_logic := 'U';
          sample_f0_35          : in    std_logic := 'U';
          sample_f0_36          : in    std_logic := 'U';
          sample_f0_37          : in    std_logic := 'U';
          sample_f0_38          : in    std_logic := 'U';
          sample_f0_39          : in    std_logic := 'U';
          sample_f0_40          : in    std_logic := 'U';
          sample_f0_41          : in    std_logic := 'U';
          sample_f0_42          : in    std_logic := 'U';
          sample_f0_43          : in    std_logic := 'U';
          sample_f0_44          : in    std_logic := 'U';
          sample_f0_45          : in    std_logic := 'U';
          sample_f0_46          : in    std_logic := 'U';
          sample_f0_47          : in    std_logic := 'U';
          sample_f0_48          : in    std_logic := 'U';
          sample_f0_49          : in    std_logic := 'U';
          sample_f0_50          : in    std_logic := 'U';
          sample_f0_51          : in    std_logic := 'U';
          sample_f0_52          : in    std_logic := 'U';
          sample_f0_53          : in    std_logic := 'U';
          sample_f0_54          : in    std_logic := 'U';
          sample_f0_55          : in    std_logic := 'U';
          sample_f0_56          : in    std_logic := 'U';
          sample_f0_57          : in    std_logic := 'U';
          sample_f0_58          : in    std_logic := 'U';
          sample_f0_59          : in    std_logic := 'U';
          sample_f0_60          : in    std_logic := 'U';
          sample_f0_61          : in    std_logic := 'U';
          sample_f0_62          : in    std_logic := 'U';
          sample_f0_63          : in    std_logic := 'U';
          sample_f1_0           : out   std_logic;
          sample_f1_1           : out   std_logic;
          sample_f1_2           : out   std_logic;
          sample_f1_3           : out   std_logic;
          sample_f1_4           : out   std_logic;
          sample_f1_5           : out   std_logic;
          sample_f1_6           : out   std_logic;
          sample_f1_7           : out   std_logic;
          sample_f1_8           : out   std_logic;
          sample_f1_9           : out   std_logic;
          sample_f1_10          : out   std_logic;
          sample_f1_11          : out   std_logic;
          sample_f1_12          : out   std_logic;
          sample_f1_13          : out   std_logic;
          sample_f1_14          : out   std_logic;
          sample_f1_15          : out   std_logic;
          sample_f1_32          : out   std_logic;
          sample_f1_33          : out   std_logic;
          sample_f1_34          : out   std_logic;
          sample_f1_35          : out   std_logic;
          sample_f1_36          : out   std_logic;
          sample_f1_37          : out   std_logic;
          sample_f1_38          : out   std_logic;
          sample_f1_39          : out   std_logic;
          sample_f1_40          : out   std_logic;
          sample_f1_41          : out   std_logic;
          sample_f1_42          : out   std_logic;
          sample_f1_43          : out   std_logic;
          sample_f1_44          : out   std_logic;
          sample_f1_45          : out   std_logic;
          sample_f1_46          : out   std_logic;
          sample_f1_47          : out   std_logic;
          sample_f1_48          : out   std_logic;
          sample_f1_49          : out   std_logic;
          sample_f1_50          : out   std_logic;
          sample_f1_51          : out   std_logic;
          sample_f1_52          : out   std_logic;
          sample_f1_53          : out   std_logic;
          sample_f1_54          : out   std_logic;
          sample_f1_55          : out   std_logic;
          sample_f1_56          : out   std_logic;
          sample_f1_57          : out   std_logic;
          sample_f1_58          : out   std_logic;
          sample_f1_59          : out   std_logic;
          sample_f1_60          : out   std_logic;
          sample_f1_61          : out   std_logic;
          sample_f1_62          : out   std_logic;
          sample_f1_63          : out   std_logic;
          sample_f0_wdata_95    : in    std_logic := 'U';
          sample_f0_wdata_94    : in    std_logic := 'U';
          sample_f0_wdata_93    : in    std_logic := 'U';
          sample_f0_wdata_92    : in    std_logic := 'U';
          sample_f0_wdata_91    : in    std_logic := 'U';
          sample_f0_wdata_90    : in    std_logic := 'U';
          sample_f0_wdata_89    : in    std_logic := 'U';
          sample_f0_wdata_88    : in    std_logic := 'U';
          sample_f0_wdata_87    : in    std_logic := 'U';
          sample_f0_wdata_86    : in    std_logic := 'U';
          sample_f0_wdata_85    : in    std_logic := 'U';
          sample_f0_wdata_84    : in    std_logic := 'U';
          sample_f0_wdata_83    : in    std_logic := 'U';
          sample_f0_wdata_82    : in    std_logic := 'U';
          sample_f0_wdata_81    : in    std_logic := 'U';
          sample_f0_wdata_80    : in    std_logic := 'U';
          sample_f0_wdata_79    : in    std_logic := 'U';
          sample_f0_wdata_78    : in    std_logic := 'U';
          sample_f0_wdata_77    : in    std_logic := 'U';
          sample_f0_wdata_76    : in    std_logic := 'U';
          sample_f0_wdata_75    : in    std_logic := 'U';
          sample_f0_wdata_74    : in    std_logic := 'U';
          sample_f0_wdata_73    : in    std_logic := 'U';
          sample_f0_wdata_72    : in    std_logic := 'U';
          sample_f0_wdata_71    : in    std_logic := 'U';
          sample_f0_wdata_70    : in    std_logic := 'U';
          sample_f0_wdata_69    : in    std_logic := 'U';
          sample_f0_wdata_68    : in    std_logic := 'U';
          sample_f0_wdata_67    : in    std_logic := 'U';
          sample_f0_wdata_66    : in    std_logic := 'U';
          sample_f0_wdata_65    : in    std_logic := 'U';
          sample_f0_wdata_64    : in    std_logic := 'U';
          sample_f0_wdata_63    : in    std_logic := 'U';
          sample_f0_wdata_62    : in    std_logic := 'U';
          sample_f0_wdata_61    : in    std_logic := 'U';
          sample_f0_wdata_60    : in    std_logic := 'U';
          sample_f0_wdata_59    : in    std_logic := 'U';
          sample_f0_wdata_58    : in    std_logic := 'U';
          sample_f0_wdata_57    : in    std_logic := 'U';
          sample_f0_wdata_56    : in    std_logic := 'U';
          sample_f0_wdata_55    : in    std_logic := 'U';
          sample_f0_wdata_54    : in    std_logic := 'U';
          sample_f0_wdata_53    : in    std_logic := 'U';
          sample_f0_wdata_52    : in    std_logic := 'U';
          sample_f0_wdata_51    : in    std_logic := 'U';
          sample_f0_wdata_50    : in    std_logic := 'U';
          sample_f0_wdata_49    : in    std_logic := 'U';
          sample_f0_wdata_48    : in    std_logic := 'U';
          sample_f0_wdata_15    : in    std_logic := 'U';
          sample_f0_wdata_14    : in    std_logic := 'U';
          sample_f0_wdata_13    : in    std_logic := 'U';
          sample_f0_wdata_12    : in    std_logic := 'U';
          sample_f0_wdata_11    : in    std_logic := 'U';
          sample_f0_wdata_10    : in    std_logic := 'U';
          sample_f0_wdata_9     : in    std_logic := 'U';
          sample_f0_wdata_8     : in    std_logic := 'U';
          sample_f0_wdata_7     : in    std_logic := 'U';
          sample_f0_wdata_6     : in    std_logic := 'U';
          sample_f0_wdata_5     : in    std_logic := 'U';
          sample_f0_wdata_4     : in    std_logic := 'U';
          sample_f0_wdata_3     : in    std_logic := 'U';
          sample_f0_wdata_2     : in    std_logic := 'U';
          sample_f0_wdata_1     : in    std_logic := 'U';
          sample_f0_wdata_0     : in    std_logic := 'U';
          sample_f1_wdata_95    : out   std_logic;
          sample_f1_wdata_94    : out   std_logic;
          sample_f1_wdata_93    : out   std_logic;
          sample_f1_wdata_92    : out   std_logic;
          sample_f1_wdata_91    : out   std_logic;
          sample_f1_wdata_90    : out   std_logic;
          sample_f1_wdata_89    : out   std_logic;
          sample_f1_wdata_88    : out   std_logic;
          sample_f1_wdata_87    : out   std_logic;
          sample_f1_wdata_86    : out   std_logic;
          sample_f1_wdata_85    : out   std_logic;
          sample_f1_wdata_84    : out   std_logic;
          sample_f1_wdata_83    : out   std_logic;
          sample_f1_wdata_82    : out   std_logic;
          sample_f1_wdata_81    : out   std_logic;
          sample_f1_wdata_80    : out   std_logic;
          sample_f1_wdata_79    : out   std_logic;
          sample_f1_wdata_78    : out   std_logic;
          sample_f1_wdata_77    : out   std_logic;
          sample_f1_wdata_76    : out   std_logic;
          sample_f1_wdata_75    : out   std_logic;
          sample_f1_wdata_74    : out   std_logic;
          sample_f1_wdata_73    : out   std_logic;
          sample_f1_wdata_72    : out   std_logic;
          sample_f1_wdata_71    : out   std_logic;
          sample_f1_wdata_70    : out   std_logic;
          sample_f1_wdata_69    : out   std_logic;
          sample_f1_wdata_68    : out   std_logic;
          sample_f1_wdata_67    : out   std_logic;
          sample_f1_wdata_66    : out   std_logic;
          sample_f1_wdata_65    : out   std_logic;
          sample_f1_wdata_64    : out   std_logic;
          sample_f1_wdata_63    : out   std_logic;
          sample_f1_wdata_62    : out   std_logic;
          sample_f1_wdata_61    : out   std_logic;
          sample_f1_wdata_60    : out   std_logic;
          sample_f1_wdata_59    : out   std_logic;
          sample_f1_wdata_58    : out   std_logic;
          sample_f1_wdata_57    : out   std_logic;
          sample_f1_wdata_56    : out   std_logic;
          sample_f1_wdata_55    : out   std_logic;
          sample_f1_wdata_54    : out   std_logic;
          sample_f1_wdata_53    : out   std_logic;
          sample_f1_wdata_52    : out   std_logic;
          sample_f1_wdata_51    : out   std_logic;
          sample_f1_wdata_50    : out   std_logic;
          sample_f1_wdata_49    : out   std_logic;
          sample_f1_wdata_48    : out   std_logic;
          sample_f1_wdata_15    : out   std_logic;
          sample_f1_wdata_14    : out   std_logic;
          sample_f1_wdata_13    : out   std_logic;
          sample_f1_wdata_12    : out   std_logic;
          sample_f1_wdata_11    : out   std_logic;
          sample_f1_wdata_10    : out   std_logic;
          sample_f1_wdata_9     : out   std_logic;
          sample_f1_wdata_8     : out   std_logic;
          sample_f1_wdata_7     : out   std_logic;
          sample_f1_wdata_6     : out   std_logic;
          sample_f1_wdata_5     : out   std_logic;
          sample_f1_wdata_4     : out   std_logic;
          sample_f1_wdata_3     : out   std_logic;
          sample_f1_wdata_2     : out   std_logic;
          sample_f1_wdata_1     : out   std_logic;
          sample_f1_wdata_0     : out   std_logic;
          sample_f0_val_1       : in    std_logic := 'U';
          sample_f1_val         : out   std_logic;
          sample_f0_val_0       : in    std_logic := 'U';
          sample_out_0_sqmuxa_1 : out   std_logic;
          HRESETn_c             : in    std_logic := 'U';
          HCLK_c                : in    std_logic := 'U';
          sample_f1_val_0       : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AD7688_drvr
    port( sample_7   : out   std_logic_vector(15 downto 0);
          sample_0   : out   std_logic_vector(15 downto 0);
          sample_1   : out   std_logic_vector(15 downto 0);
          sample_2   : out   std_logic_vector(15 downto 0);
          sample_3   : out   std_logic_vector(15 downto 0);
          sample_4   : out   std_logic_vector(15 downto 0);
          sample_5   : out   std_logic_vector(15 downto 0);
          sdo_c      : in    std_logic_vector(7 downto 0) := (others => 'U');
          sample_6   : out   std_logic_vector(15 downto 0);
          cnv_rstn_c : in    std_logic := 'U';
          cnv_clk_c  : in    std_logic := 'U';
          cnv_c      : out   std_logic;
          sample_val : out   std_logic;
          sck_c      : out   std_logic;
          cnv_run_c  : in    std_logic := 'U';
          HRESETn_c  : in    std_logic := 'U';
          HCLK_c     : in    std_logic := 'U'
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sample_data_shaping_out_val_0\, 
        sample_filter_v2_out_val, \sample_val_delay\, 
        sample_val_delay_0, SUB_16x16_medium_area_I57_Y_2, N244, 
        N229, SUB_16x16_medium_area_I57_Y_1, N254, N212, 
        SUB_16x16_medium_area_I57_Y_0, N206, 
        \sample_filter_v2_out[111]\, \sample_filter_v2_out[93]\, 
        SUB_16x16_medium_area_I57_Y_2_0, N244_0, N229_0, 
        SUB_16x16_medium_area_I57_Y_1_0, N212_0, N254_0, 
        SUB_16x16_medium_area_I57_Y_0_0, N206_0, 
        \sample_filter_v2_out[129]\, 
        SUB_16x16_medium_area_I57_un1_Y_0, N245, 
        SUB_16x16_medium_area_I57_un1_Y_0_0, N245_0, 
        SUB_16x16_medium_area_I56_Y_1, N274, N220, 
        SUB_16x16_medium_area_I56_Y_0, N190, 
        \sample_filter_v2_out[119]\, \sample_filter_v2_out[101]\, 
        SUB_16x16_medium_area_I56_Y_1_0, N274_0, N220_0, 
        SUB_16x16_medium_area_I56_Y_0_0, N190_0, 
        \sample_filter_v2_out[137]\, 
        SUB_16x16_medium_area_I56_un1_Y_0, N275, 
        SUB_16x16_medium_area_I49_Y_0, N198, 
        \sample_filter_v2_out[115]\, \sample_filter_v2_out[97]\, 
        SUB_16x16_medium_area_I49_Y_0_0, N198_0, 
        \sample_filter_v2_out[133]\, 
        SUB_16x16_medium_area_I53_Y_0, N182, 
        \sample_filter_v2_out[123]\, \sample_filter_v2_out[105]\, 
        SUB_16x16_medium_area_I53_Y_0_0, N182_0, 
        \sample_filter_v2_out[141]\, 
        SUB_16x16_medium_area_I53_un1_Y_0, N225, N264, N216, N240, 
        N268, I53_un1_Y, N225_0, N183, N181, N278, N264_0, N216_0, 
        N240_0, N268_0, I56_un1_Y, N275_0, N278_0, 
        \sample_data_shaping_f2_f1_s[15]\, 
        \sample_filter_v2_out[110]\, \sample_filter_v2_out[92]\, 
        \sample_data_shaping_f1_f0_s[15]\, 
        \sample_filter_v2_out[128]\, N181_0, N194, 
        \sample_filter_v2_out[118]\, \sample_filter_v2_out[136]\, 
        \sample_filter_v2_out[116]\, \sample_filter_v2_out[134]\, 
        N202, \sample_filter_v2_out[114]\, 
        \sample_filter_v2_out[132]\, \sample_filter_v2_out[112]\, 
        \sample_filter_v2_out[130]\, N205, 
        \sample_filter_v2_out[131]\, \sample_filter_v2_out[113]\, 
        N255, N201, N197, N265, N195, N258, N260, N270, N282_i, 
        N284_i, N286_i, \sample_data_shaping_f1_f0_s[7]\, 
        \sample_data_shaping_f1_f0_s[9]\, 
        \sample_data_shaping_f1_f0_s[10]\, 
        \sample_data_shaping_f1_f0_s[11]\, 
        \sample_data_shaping_f1_f0_s[12]\, 
        \sample_data_shaping_f1_f0_s[13]\, 
        \sample_data_shaping_f1_f0_s_i[14]\, N186, 
        \sample_filter_v2_out[122]\, \sample_filter_v2_out[140]\, 
        \sample_filter_v2_out[120]\, \sample_filter_v2_out[138]\, 
        N191, N189, \sample_filter_v2_out[121]\, 
        \sample_filter_v2_out[139]\, N187, N185, I85_un1_Y, 
        I90_un1_Y, SUB_16x16_medium_area_I91_un1_Y, 
        \sample_data_shaping_f1_f0_s[3]\, 
        \sample_data_shaping_f1_f0_s[4]\, 
        \sample_data_shaping_f1_f0_s[5]\, 
        \sample_data_shaping_f1_f0_s[6]\, N194_0, 
        \sample_filter_v2_out[100]\, \sample_filter_v2_out[98]\, 
        N202_0, \sample_filter_v2_out[96]\, 
        \sample_filter_v2_out[94]\, N207, N205_0, 
        \sample_filter_v2_out[95]\, N255_0, N203, N201_0, N199, 
        N197_0, \sample_filter_v2_out[99]\, 
        \sample_filter_v2_out[117]\, N265_0, N195_0, N193, 
        I64_un1_Y, I71_un1_Y, I78_un1_Y, I86_un1_Y, 
        SUB_16x16_medium_area_I87_un1_Y, I88_un1_Y, 
        SUB_16x16_medium_area_I89_un1_Y, 
        \sample_data_shaping_f2_f1_s[7]\, 
        \sample_data_shaping_f2_f1_s[8]\, 
        \sample_data_shaping_f2_f1_s[9]\, 
        \sample_data_shaping_f2_f1_s[10]\, 
        \sample_data_shaping_f2_f1_s[11]\, 
        \sample_data_shaping_f2_f1_s[12]\, 
        \sample_data_shaping_f2_f1_s[13]\, 
        \sample_data_shaping_f2_f1_s[14]\, N186_0, 
        \sample_filter_v2_out[104]\, \sample_filter_v2_out[102]\, 
        N189_0, \sample_filter_v2_out[103]\, N187_0, N280, N290_i, 
        SUB_16x16_medium_area_I91_un1_Y_0, 
        \sample_data_shaping_f2_f1_s[3]\, 
        \sample_data_shaping_f2_f1_s[4]\, 
        \sample_data_shaping_f2_f1_s[5]\, 
        \sample_data_shaping_f2_f1_s[6]\, 
        \sample_data_shaping_out_377[92]\, 
        \sample_data_shaping_out_353[93]\, 
        \sample_data_shaping_out_329[94]\, 
        \sample_data_shaping_out_305[95]\, 
        \sample_data_shaping_out_281[96]\, 
        \sample_data_shaping_out_257[97]\, 
        \sample_data_shaping_out_233[98]\, 
        \sample_data_shaping_out_209[99]\, 
        \sample_data_shaping_out_185[100]\, 
        \sample_data_shaping_out_161[101]\, 
        \sample_data_shaping_out_137[102]\, 
        \sample_data_shaping_out_113[103]\, 
        \sample_data_shaping_out_89[104]\, 
        \sample_data_shaping_out_373[110]\, 
        \sample_data_shaping_out_349[111]\, 
        \sample_data_shaping_out_325[112]\, 
        \sample_data_shaping_out_301[113]\, 
        \sample_data_shaping_out_277[114]\, 
        \sample_data_shaping_out_253[115]\, 
        \sample_data_shaping_out_229[116]\, 
        \sample_data_shaping_out_181[118]\, 
        \sample_data_shaping_out_157[119]\, 
        \sample_data_shaping_out_133[120]\, 
        \sample_data_shaping_out_109[121]\, 
        \sample_data_shaping_out_85[122]\, 
        \sample_filter_v2_out[143]\, \sample_filter_v2_out[125]\, 
        \sample_filter_v2_out[107]\, 
        \sample_data_shaping_out_17[107]\, 
        \sample_data_shaping_out_13[125]\, 
        \sample_data_shaping_out_37[124]\, 
        \sample_filter_v2_out[124]\, 
        \sample_data_shaping_f1_f0_s[1]\, 
        \sample_data_shaping_out_61[123]\, 
        \sample_data_shaping_f1_f0_s[2]\, 
        \sample_data_shaping_out_205[117]\, 
        \sample_data_shaping_f1_f0_s[8]\, 
        \sample_data_shaping_out_41[106]\, 
        \sample_filter_v2_out[106]\, 
        \sample_data_shaping_f2_f1_s[1]\, 
        \sample_data_shaping_out_65[105]\, 
        \sample_data_shaping_f2_f1_s[2]\, N294_i, I92_un1_Y, 
        \sample_filter_v2_out[142]\, \sample_filter_v2_out[135]\, 
        N288_i, sample_val, \sample_data_shaping_out_val\, 
        \sample_data_shaping_out[20]\, \sample_filter_v2_out[20]\, 
        \sample_data_shaping_out[21]\, \sample_filter_v2_out[21]\, 
        \sample_data_shaping_out[22]\, \sample_filter_v2_out[22]\, 
        \sample_data_shaping_out[23]\, \sample_filter_v2_out[23]\, 
        \sample_data_shaping_out[24]\, \sample_filter_v2_out[24]\, 
        \sample_data_shaping_out[25]\, \sample_filter_v2_out[25]\, 
        \sample_data_shaping_out[26]\, \sample_filter_v2_out[26]\, 
        \sample_data_shaping_out[27]\, \sample_filter_v2_out[27]\, 
        \sample_data_shaping_out[28]\, \sample_filter_v2_out[28]\, 
        \sample_data_shaping_out[29]\, \sample_filter_v2_out[29]\, 
        \sample_data_shaping_out[30]\, \sample_filter_v2_out[30]\, 
        \sample_data_shaping_out[31]\, \sample_filter_v2_out[31]\, 
        \sample_data_shaping_out[32]\, \sample_filter_v2_out[32]\, 
        \sample_data_shaping_out[33]\, \sample_filter_v2_out[33]\, 
        \sample_data_shaping_out[34]\, \sample_filter_v2_out[34]\, 
        \sample_data_shaping_out[35]\, \sample_filter_v2_out[35]\, 
        \sample_data_shaping_out[38]\, \sample_filter_v2_out[38]\, 
        \sample_data_shaping_out[39]\, \sample_filter_v2_out[39]\, 
        \sample_data_shaping_out[40]\, \sample_filter_v2_out[40]\, 
        \sample_data_shaping_out[41]\, \sample_filter_v2_out[41]\, 
        \sample_data_shaping_out[42]\, \sample_filter_v2_out[42]\, 
        \sample_data_shaping_out[43]\, \sample_filter_v2_out[43]\, 
        \sample_data_shaping_out[44]\, \sample_filter_v2_out[44]\, 
        \sample_data_shaping_out[45]\, \sample_filter_v2_out[45]\, 
        \sample_data_shaping_out[46]\, \sample_filter_v2_out[46]\, 
        \sample_data_shaping_out[47]\, \sample_filter_v2_out[47]\, 
        \sample_data_shaping_out[48]\, \sample_filter_v2_out[48]\, 
        \sample_data_shaping_out[49]\, \sample_filter_v2_out[49]\, 
        \sample_data_shaping_out[50]\, \sample_filter_v2_out[50]\, 
        \sample_data_shaping_out[51]\, \sample_filter_v2_out[51]\, 
        \sample_data_shaping_out[52]\, \sample_filter_v2_out[52]\, 
        \sample_data_shaping_out[53]\, \sample_filter_v2_out[53]\, 
        \sample_data_shaping_out[56]\, \sample_filter_v2_out[56]\, 
        \sample_data_shaping_out[57]\, \sample_filter_v2_out[57]\, 
        \sample_data_shaping_out[58]\, \sample_filter_v2_out[58]\, 
        \sample_data_shaping_out[59]\, \sample_filter_v2_out[59]\, 
        \sample_data_shaping_out[60]\, \sample_filter_v2_out[60]\, 
        \sample_data_shaping_out[61]\, \sample_filter_v2_out[61]\, 
        \sample_data_shaping_out[62]\, \sample_filter_v2_out[62]\, 
        \sample_data_shaping_out[63]\, \sample_filter_v2_out[63]\, 
        \sample_data_shaping_out[64]\, \sample_filter_v2_out[64]\, 
        \sample_data_shaping_out[65]\, \sample_filter_v2_out[65]\, 
        \sample_data_shaping_out[66]\, \sample_filter_v2_out[66]\, 
        \sample_data_shaping_out[67]\, \sample_filter_v2_out[67]\, 
        \sample_data_shaping_out[68]\, \sample_filter_v2_out[68]\, 
        \sample_data_shaping_out[69]\, \sample_filter_v2_out[69]\, 
        \sample_data_shaping_out[70]\, \sample_filter_v2_out[70]\, 
        \sample_data_shaping_out[71]\, \sample_filter_v2_out[71]\, 
        \sample_data_shaping_out[128]\, 
        \sample_data_shaping_out[129]\, 
        \sample_data_shaping_out[130]\, 
        \sample_data_shaping_out[131]\, 
        \sample_data_shaping_out[132]\, 
        \sample_data_shaping_out[133]\, 
        \sample_data_shaping_out[134]\, 
        \sample_data_shaping_out[135]\, 
        \sample_data_shaping_out[136]\, 
        \sample_data_shaping_out[137]\, 
        \sample_data_shaping_out[138]\, 
        \sample_data_shaping_out[139]\, 
        \sample_data_shaping_out[140]\, 
        \sample_data_shaping_out[141]\, 
        \sample_data_shaping_out[142]\, 
        \sample_data_shaping_out[143]\, 
        \sample_data_shaping_out[2]\, \sample_filter_v2_out[2]\, 
        \sample_data_shaping_out[3]\, \sample_filter_v2_out[3]\, 
        \sample_data_shaping_out[4]\, \sample_filter_v2_out[4]\, 
        \sample_data_shaping_out[5]\, \sample_filter_v2_out[5]\, 
        \sample_data_shaping_out[6]\, \sample_filter_v2_out[6]\, 
        \sample_data_shaping_out[7]\, \sample_filter_v2_out[7]\, 
        \sample_data_shaping_out[8]\, \sample_filter_v2_out[8]\, 
        \sample_data_shaping_out[9]\, \sample_filter_v2_out[9]\, 
        \sample_data_shaping_out[10]\, \sample_filter_v2_out[10]\, 
        \sample_data_shaping_out[11]\, \sample_filter_v2_out[11]\, 
        \sample_data_shaping_out[12]\, \sample_filter_v2_out[12]\, 
        \sample_data_shaping_out[13]\, \sample_filter_v2_out[13]\, 
        \sample_data_shaping_out[14]\, \sample_filter_v2_out[14]\, 
        \sample_data_shaping_out[15]\, \sample_filter_v2_out[15]\, 
        \sample_data_shaping_out[16]\, \sample_filter_v2_out[16]\, 
        \sample_data_shaping_out[17]\, \sample_filter_v2_out[17]\, 
        \sample_data_shaping_out[92]\, 
        \sample_data_shaping_out[93]\, 
        \sample_data_shaping_out[94]\, 
        \sample_data_shaping_out[95]\, 
        \sample_data_shaping_out[96]\, 
        \sample_data_shaping_out[97]\, 
        \sample_data_shaping_out[98]\, 
        \sample_data_shaping_out[99]\, 
        \sample_data_shaping_out[100]\, 
        \sample_data_shaping_out[101]\, 
        \sample_data_shaping_out[102]\, 
        \sample_data_shaping_out[103]\, 
        \sample_data_shaping_out[104]\, 
        \sample_data_shaping_out[105]\, 
        \sample_data_shaping_out[106]\, 
        \sample_data_shaping_out[107]\, 
        \sample_data_shaping_out[110]\, 
        \sample_data_shaping_out[111]\, 
        \sample_data_shaping_out[112]\, 
        \sample_data_shaping_out[113]\, 
        \sample_data_shaping_out[114]\, 
        \sample_data_shaping_out[115]\, 
        \sample_data_shaping_out[116]\, 
        \sample_data_shaping_out[117]\, 
        \sample_data_shaping_out[118]\, 
        \sample_data_shaping_out[119]\, 
        \sample_data_shaping_out[120]\, 
        \sample_data_shaping_out[121]\, 
        \sample_data_shaping_out[122]\, 
        \sample_data_shaping_out[123]\, 
        \sample_data_shaping_out[124]\, 
        \sample_data_shaping_out[125]\, \sample_7[0]\, 
        \sample_7[1]\, \sample_7[2]\, \sample_7[3]\, 
        \sample_7[4]\, \sample_7[5]\, \sample_7[6]\, 
        \sample_7[7]\, \sample_7[8]\, \sample_7[9]\, 
        \sample_7[10]\, \sample_7[11]\, \sample_7[12]\, 
        \sample_7[13]\, \sample_7[14]\, \sample_7[15]\, 
        \sample_0[0]\, \sample_0[1]\, \sample_0[2]\, 
        \sample_0[3]\, \sample_0[4]\, \sample_0[5]\, 
        \sample_0[6]\, \sample_0[7]\, \sample_0[8]\, 
        \sample_0[9]\, \sample_0[10]\, \sample_0[11]\, 
        \sample_0[12]\, \sample_0[13]\, \sample_0[14]\, 
        \sample_0[15]\, \sample_1[0]\, \sample_1[1]\, 
        \sample_1[2]\, \sample_1[3]\, \sample_1[4]\, 
        \sample_1[5]\, \sample_1[6]\, \sample_1[7]\, 
        \sample_1[8]\, \sample_1[9]\, \sample_1[10]\, 
        \sample_1[11]\, \sample_1[12]\, \sample_1[13]\, 
        \sample_1[14]\, \sample_1[15]\, \sample_2[0]\, 
        \sample_2[1]\, \sample_2[2]\, \sample_2[3]\, 
        \sample_2[4]\, \sample_2[5]\, \sample_2[6]\, 
        \sample_2[7]\, \sample_2[8]\, \sample_2[9]\, 
        \sample_2[10]\, \sample_2[11]\, \sample_2[12]\, 
        \sample_2[13]\, \sample_2[14]\, \sample_2[15]\, 
        \sample_3[0]\, \sample_3[1]\, \sample_3[2]\, 
        \sample_3[3]\, \sample_3[4]\, \sample_3[5]\, 
        \sample_3[6]\, \sample_3[7]\, \sample_3[8]\, 
        \sample_3[9]\, \sample_3[10]\, \sample_3[11]\, 
        \sample_3[12]\, \sample_3[13]\, \sample_3[14]\, 
        \sample_3[15]\, \sample_4[0]\, \sample_4[1]\, 
        \sample_4[2]\, \sample_4[3]\, \sample_4[4]\, 
        \sample_4[5]\, \sample_4[6]\, \sample_4[7]\, 
        \sample_4[8]\, \sample_4[9]\, \sample_4[10]\, 
        \sample_4[11]\, \sample_4[12]\, \sample_4[13]\, 
        \sample_4[14]\, \sample_4[15]\, \sample_5[0]\, 
        \sample_5[1]\, \sample_5[2]\, \sample_5[3]\, 
        \sample_5[4]\, \sample_5[5]\, \sample_5[6]\, 
        \sample_5[7]\, \sample_5[8]\, \sample_5[9]\, 
        \sample_5[10]\, \sample_5[11]\, \sample_5[12]\, 
        \sample_5[13]\, \sample_5[14]\, \sample_5[15]\, 
        \sample_6[0]\, \sample_6[1]\, \sample_6[2]\, 
        \sample_6[3]\, \sample_6[4]\, \sample_6[5]\, 
        \sample_6[6]\, \sample_6[7]\, \sample_6[8]\, 
        \sample_6[9]\, \sample_6[10]\, \sample_6[11]\, 
        \sample_6[12]\, \sample_6[13]\, \sample_6[14]\, 
        \sample_6[15]\, \sample_f0[48]\, \sample_f0[49]\, 
        \sample_f0[50]\, \sample_f0[51]\, \sample_f0[52]\, 
        \sample_f0[53]\, \sample_f0[54]\, \sample_f0[55]\, 
        \sample_f0[56]\, \sample_f0[57]\, \sample_f0[58]\, 
        \sample_f0[59]\, \sample_f0[60]\, \sample_f0[61]\, 
        \sample_f0[62]\, \sample_f0[63]\, \sample_f0[80]\, 
        \sample_f0[81]\, \sample_f0[82]\, \sample_f0[83]\, 
        \sample_f0[84]\, \sample_f0[85]\, \sample_f0[86]\, 
        \sample_f0[87]\, \sample_f0[88]\, \sample_f0[89]\, 
        \sample_f0[90]\, \sample_f0[91]\, \sample_f0[92]\, 
        \sample_f0[93]\, \sample_f0[94]\, \sample_f0[95]\, 
        \sample_f0[96]\, \sample_f0[97]\, \sample_f0[98]\, 
        \sample_f0[99]\, \sample_f0[100]\, \sample_f0[101]\, 
        \sample_f0[102]\, \sample_f0[103]\, \sample_f0[104]\, 
        \sample_f0[105]\, \sample_f0[106]\, \sample_f0[107]\, 
        \sample_f0[108]\, \sample_f0[109]\, \sample_f0[110]\, 
        \sample_f0[111]\, \sample_f0_wdata[95]\, 
        \sample_f0_wdata[94]\, \sample_f0_wdata[93]\, 
        \sample_f0_wdata[92]\, \sample_f0_wdata[91]\, 
        \sample_f0_wdata[90]\, \sample_f0_wdata[89]\, 
        \sample_f0_wdata[88]\, \sample_f0_wdata[87]\, 
        \sample_f0_wdata[86]\, \sample_f0_wdata[85]\, 
        \sample_f0_wdata[84]\, \sample_f0_wdata[83]\, 
        \sample_f0_wdata[82]\, \sample_f0_wdata[81]\, 
        \sample_f0_wdata[80]\, \sample_f0_wdata[79]\, 
        \sample_f0_wdata[78]\, \sample_f0_wdata[77]\, 
        \sample_f0_wdata[76]\, \sample_f0_wdata[75]\, 
        \sample_f0_wdata[74]\, \sample_f0_wdata[73]\, 
        \sample_f0_wdata[72]\, \sample_f0_wdata[71]\, 
        \sample_f0_wdata[70]\, \sample_f0_wdata[69]\, 
        \sample_f0_wdata[68]\, \sample_f0_wdata[67]\, 
        \sample_f0_wdata[66]\, \sample_f0_wdata[65]\, 
        \sample_f0_wdata[64]\, \sample_f0_wdata[63]\, 
        \sample_f0_wdata[62]\, \sample_f0_wdata[61]\, 
        \sample_f0_wdata[60]\, \sample_f0_wdata[59]\, 
        \sample_f0_wdata[58]\, \sample_f0_wdata[57]\, 
        \sample_f0_wdata[56]\, \sample_f0_wdata[55]\, 
        \sample_f0_wdata[54]\, \sample_f0_wdata[53]\, 
        \sample_f0_wdata[52]\, \sample_f0_wdata[51]\, 
        \sample_f0_wdata[50]\, \sample_f0_wdata[49]\, 
        \sample_f0_wdata[48]\, \sample_f0_wdata[15]\, 
        \sample_f0_wdata[14]\, \sample_f0_wdata[13]\, 
        \sample_f0_wdata[12]\, \sample_f0_wdata[11]\, 
        \sample_f0_wdata[10]\, \sample_f0_wdata[9]\, 
        \sample_f0_wdata[8]\, \sample_f0_wdata[7]\, 
        \sample_f0_wdata[6]\, \sample_f0_wdata[5]\, 
        \sample_f0_wdata[4]\, \sample_f0_wdata[3]\, 
        \sample_f0_wdata[2]\, \sample_f0_wdata[1]\, 
        \sample_f0_wdata[0]\, sample_f0_val, sample_f0_val_0, 
        sample_f0_val_1, \sample_f1[48]\, \sample_f1[49]\, 
        \sample_f1[50]\, \sample_f1[51]\, \sample_f1[52]\, 
        \sample_f1[53]\, \sample_f1[54]\, \sample_f1[55]\, 
        \sample_f1[56]\, \sample_f1[57]\, \sample_f1[58]\, 
        \sample_f1[59]\, \sample_f1[60]\, \sample_f1[61]\, 
        \sample_f1[62]\, \sample_f1[63]\, \sample_f1[80]\, 
        \sample_f1[81]\, \sample_f1[82]\, \sample_f1[83]\, 
        \sample_f1[84]\, \sample_f1[85]\, \sample_f1[86]\, 
        \sample_f1[87]\, \sample_f1[88]\, \sample_f1[89]\, 
        \sample_f1[90]\, \sample_f1[91]\, \sample_f1[92]\, 
        \sample_f1[93]\, \sample_f1[94]\, \sample_f1[95]\, 
        \sample_f1[96]\, \sample_f1[97]\, \sample_f1[98]\, 
        \sample_f1[99]\, \sample_f1[100]\, \sample_f1[101]\, 
        \sample_f1[102]\, \sample_f1[103]\, \sample_f1[104]\, 
        \sample_f1[105]\, \sample_f1[106]\, \sample_f1[107]\, 
        \sample_f1[108]\, \sample_f1[109]\, \sample_f1[110]\, 
        \sample_f1[111]\, \sample_f1_wdata[95]\, 
        \sample_f1_wdata[94]\, \sample_f1_wdata[93]\, 
        \sample_f1_wdata[92]\, \sample_f1_wdata[91]\, 
        \sample_f1_wdata[90]\, \sample_f1_wdata[89]\, 
        \sample_f1_wdata[88]\, \sample_f1_wdata[87]\, 
        \sample_f1_wdata[86]\, \sample_f1_wdata[85]\, 
        \sample_f1_wdata[84]\, \sample_f1_wdata[83]\, 
        \sample_f1_wdata[82]\, \sample_f1_wdata[81]\, 
        \sample_f1_wdata[80]\, \sample_f1_wdata[79]\, 
        \sample_f1_wdata[78]\, \sample_f1_wdata[77]\, 
        \sample_f1_wdata[76]\, \sample_f1_wdata[75]\, 
        \sample_f1_wdata[74]\, \sample_f1_wdata[73]\, 
        \sample_f1_wdata[72]\, \sample_f1_wdata[71]\, 
        \sample_f1_wdata[70]\, \sample_f1_wdata[69]\, 
        \sample_f1_wdata[68]\, \sample_f1_wdata[67]\, 
        \sample_f1_wdata[66]\, \sample_f1_wdata[65]\, 
        \sample_f1_wdata[64]\, \sample_f1_wdata[63]\, 
        \sample_f1_wdata[62]\, \sample_f1_wdata[61]\, 
        \sample_f1_wdata[60]\, \sample_f1_wdata[59]\, 
        \sample_f1_wdata[58]\, \sample_f1_wdata[57]\, 
        \sample_f1_wdata[56]\, \sample_f1_wdata[55]\, 
        \sample_f1_wdata[54]\, \sample_f1_wdata[53]\, 
        \sample_f1_wdata[52]\, \sample_f1_wdata[51]\, 
        \sample_f1_wdata[50]\, \sample_f1_wdata[49]\, 
        \sample_f1_wdata[48]\, \sample_f1_wdata[15]\, 
        \sample_f1_wdata[14]\, \sample_f1_wdata[13]\, 
        \sample_f1_wdata[12]\, \sample_f1_wdata[11]\, 
        \sample_f1_wdata[10]\, \sample_f1_wdata[9]\, 
        \sample_f1_wdata[8]\, \sample_f1_wdata[7]\, 
        \sample_f1_wdata[6]\, \sample_f1_wdata[5]\, 
        \sample_f1_wdata[4]\, \sample_f1_wdata[3]\, 
        \sample_f1_wdata[2]\, \sample_f1_wdata[1]\, 
        \sample_f1_wdata[0]\, sample_f1_val, 
        sample_out_0_sqmuxa_1, sample_f1_val_0, 
        \sample_f2_wdata[0]\, \sample_f2_wdata[1]\, 
        \sample_f2_wdata[2]\, \sample_f2_wdata[3]\, 
        \sample_f2_wdata[4]\, \sample_f2_wdata[5]\, 
        \sample_f2_wdata[6]\, \sample_f2_wdata[7]\, 
        \sample_f2_wdata[8]\, \sample_f2_wdata[9]\, 
        \sample_f2_wdata[10]\, \sample_f2_wdata[11]\, 
        \sample_f2_wdata[12]\, \sample_f2_wdata[13]\, 
        \sample_f2_wdata[14]\, \sample_f2_wdata[15]\, 
        \sample_f2_wdata[16]\, \sample_f2_wdata[17]\, 
        \sample_f2_wdata[18]\, \sample_f2_wdata[19]\, 
        \sample_f2_wdata[20]\, \sample_f2_wdata[21]\, 
        \sample_f2_wdata[22]\, \sample_f2_wdata[23]\, 
        \sample_f2_wdata[24]\, \sample_f2_wdata[25]\, 
        \sample_f2_wdata[26]\, \sample_f2_wdata[27]\, 
        \sample_f2_wdata[28]\, \sample_f2_wdata[29]\, 
        \sample_f2_wdata[30]\, \sample_f2_wdata[31]\, 
        \sample_f2_wdata[32]\, \sample_f2_wdata[33]\, 
        \sample_f2_wdata[34]\, \sample_f2_wdata[35]\, 
        \sample_f2_wdata[36]\, \sample_f2_wdata[37]\, 
        \sample_f2_wdata[38]\, \sample_f2_wdata[39]\, 
        \sample_f2_wdata[40]\, \sample_f2_wdata[41]\, 
        \sample_f2_wdata[42]\, \sample_f2_wdata[43]\, 
        \sample_f2_wdata[44]\, \sample_f2_wdata[45]\, 
        \sample_f2_wdata[46]\, \sample_f2_wdata[47]\, 
        \sample_f2_wdata[48]\, \sample_f2_wdata[49]\, 
        \sample_f2_wdata[50]\, \sample_f2_wdata[51]\, 
        \sample_f2_wdata[52]\, \sample_f2_wdata[53]\, 
        \sample_f2_wdata[54]\, \sample_f2_wdata[55]\, 
        \sample_f2_wdata[56]\, \sample_f2_wdata[57]\, 
        \sample_f2_wdata[58]\, \sample_f2_wdata[59]\, 
        \sample_f2_wdata[60]\, \sample_f2_wdata[61]\, 
        \sample_f2_wdata[62]\, \sample_f2_wdata[63]\, 
        \sample_f2_wdata[64]\, \sample_f2_wdata[65]\, 
        \sample_f2_wdata[66]\, \sample_f2_wdata[67]\, 
        \sample_f2_wdata[68]\, \sample_f2_wdata[69]\, 
        \sample_f2_wdata[70]\, \sample_f2_wdata[71]\, 
        \sample_f2_wdata[72]\, \sample_f2_wdata[73]\, 
        \sample_f2_wdata[74]\, \sample_f2_wdata[75]\, 
        \sample_f2_wdata[76]\, \sample_f2_wdata[77]\, 
        \sample_f2_wdata[78]\, \sample_f2_wdata[79]\, 
        \sample_f2_wdata[80]\, \sample_f2_wdata[81]\, 
        \sample_f2_wdata[82]\, \sample_f2_wdata[83]\, 
        \sample_f2_wdata[84]\, \sample_f2_wdata[85]\, 
        \sample_f2_wdata[86]\, \sample_f2_wdata[87]\, 
        \sample_f2_wdata[88]\, \sample_f2_wdata[89]\, 
        \sample_f2_wdata[90]\, \sample_f2_wdata[91]\, 
        \sample_f2_wdata[92]\, \sample_f2_wdata[93]\, 
        \sample_f2_wdata[94]\, \sample_f2_wdata[95]\, 
        sample_f2_val, \sample_f3_wdata[0]\, \sample_f3_wdata[1]\, 
        \sample_f3_wdata[2]\, \sample_f3_wdata[3]\, 
        \sample_f3_wdata[4]\, \sample_f3_wdata[5]\, 
        \sample_f3_wdata[6]\, \sample_f3_wdata[7]\, 
        \sample_f3_wdata[8]\, \sample_f3_wdata[9]\, 
        \sample_f3_wdata[10]\, \sample_f3_wdata[11]\, 
        \sample_f3_wdata[12]\, \sample_f3_wdata[13]\, 
        \sample_f3_wdata[14]\, \sample_f3_wdata[15]\, 
        \sample_f3_wdata[16]\, \sample_f3_wdata[17]\, 
        \sample_f3_wdata[18]\, \sample_f3_wdata[19]\, 
        \sample_f3_wdata[20]\, \sample_f3_wdata[21]\, 
        \sample_f3_wdata[22]\, \sample_f3_wdata[23]\, 
        \sample_f3_wdata[24]\, \sample_f3_wdata[25]\, 
        \sample_f3_wdata[26]\, \sample_f3_wdata[27]\, 
        \sample_f3_wdata[28]\, \sample_f3_wdata[29]\, 
        \sample_f3_wdata[30]\, \sample_f3_wdata[31]\, 
        \sample_f3_wdata[32]\, \sample_f3_wdata[33]\, 
        \sample_f3_wdata[34]\, \sample_f3_wdata[35]\, 
        \sample_f3_wdata[36]\, \sample_f3_wdata[37]\, 
        \sample_f3_wdata[38]\, \sample_f3_wdata[39]\, 
        \sample_f3_wdata[40]\, \sample_f3_wdata[41]\, 
        \sample_f3_wdata[42]\, \sample_f3_wdata[43]\, 
        \sample_f3_wdata[44]\, \sample_f3_wdata[45]\, 
        \sample_f3_wdata[46]\, \sample_f3_wdata[47]\, 
        \sample_f3_wdata[48]\, \sample_f3_wdata[49]\, 
        \sample_f3_wdata[50]\, \sample_f3_wdata[51]\, 
        \sample_f3_wdata[52]\, \sample_f3_wdata[53]\, 
        \sample_f3_wdata[54]\, \sample_f3_wdata[55]\, 
        \sample_f3_wdata[56]\, \sample_f3_wdata[57]\, 
        \sample_f3_wdata[58]\, \sample_f3_wdata[59]\, 
        \sample_f3_wdata[60]\, \sample_f3_wdata[61]\, 
        \sample_f3_wdata[62]\, \sample_f3_wdata[63]\, 
        \sample_f3_wdata[64]\, \sample_f3_wdata[65]\, 
        \sample_f3_wdata[66]\, \sample_f3_wdata[67]\, 
        \sample_f3_wdata[68]\, \sample_f3_wdata[69]\, 
        \sample_f3_wdata[70]\, \sample_f3_wdata[71]\, 
        \sample_f3_wdata[72]\, \sample_f3_wdata[73]\, 
        \sample_f3_wdata[74]\, \sample_f3_wdata[75]\, 
        \sample_f3_wdata[76]\, \sample_f3_wdata[77]\, 
        \sample_f3_wdata[78]\, \sample_f3_wdata[79]\, 
        \sample_f3_wdata[80]\, \sample_f3_wdata[81]\, 
        \sample_f3_wdata[82]\, \sample_f3_wdata[83]\, 
        \sample_f3_wdata[84]\, \sample_f3_wdata[85]\, 
        \sample_f3_wdata[86]\, \sample_f3_wdata[87]\, 
        \sample_f3_wdata[88]\, \sample_f3_wdata[89]\, 
        \sample_f3_wdata[90]\, \sample_f3_wdata[91]\, 
        \sample_f3_wdata[92]\, \sample_f3_wdata[93]\, 
        \sample_f3_wdata[94]\, \sample_f3_wdata[95]\, 
        sample_f3_val, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : IIR_CEL_CTRLR_v2
	Use entity work.IIR_CEL_CTRLR_v2(DEF_ARCH);
    for all : Downsampling_6_16_256
	Use entity work.Downsampling_6_16_256(DEF_ARCH);
    for all : Downsampling_6_16_96
	Use entity work.Downsampling_6_16_96(DEF_ARCH);
    for all : lpp_waveform
	Use entity work.lpp_waveform(DEF_ARCH);
    for all : Downsampling_8_16_4
	Use entity work.Downsampling_8_16_4(DEF_ARCH);
    for all : Downsampling_8_16_6
	Use entity work.Downsampling_8_16_6(DEF_ARCH);
    for all : AD7688_drvr
	Use entity work.AD7688_drvr(DEF_ARCH);
begin 


    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I91_un1_Y : 
        XA1A
      port map(A => \sample_filter_v2_out[104]\, B => 
        \sample_filter_v2_out[122]\, C => N278_0, Y => 
        SUB_16x16_medium_area_I91_un1_Y_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I27_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[96]\, B => 
        \sample_filter_v2_out[114]\, Y => N202_0);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[29]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[29]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[29]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[97]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_257[97]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[97]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out_RNO[120]\ : 
        MX2
      port map(A => \sample_filter_v2_out[120]\, B => 
        \sample_data_shaping_f1_f0_s[5]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_133[120]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[138]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[138]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[138]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I86_Y : 
        AO18
      port map(A => N260, B => \sample_filter_v2_out[130]\, C => 
        \sample_filter_v2_out[112]\, Y => N282_i);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[117]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_205[117]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[117]\);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[23]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[23]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[23]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out_RNO[103]\ : 
        MX2
      port map(A => \sample_filter_v2_out[103]\, B => 
        \sample_data_shaping_f2_f1_s[4]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_113[103]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I106_Y_0 : 
        AX1D
      port map(A => I71_un1_Y, B => N254, C => N205_0, Y => 
        \sample_data_shaping_f2_f1_s[13]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I100_Y_0 : 
        XOR2
      port map(A => N268_0, B => N193, Y => 
        \sample_data_shaping_f2_f1_s[7]\);
    
    IIR_CEL_CTRLR_v2_1 : IIR_CEL_CTRLR_v2
      port map(sample_filter_v2_out_0 => 
        \sample_filter_v2_out[2]\, sample_filter_v2_out_1 => 
        \sample_filter_v2_out[3]\, sample_filter_v2_out_2 => 
        \sample_filter_v2_out[4]\, sample_filter_v2_out_3 => 
        \sample_filter_v2_out[5]\, sample_filter_v2_out_4 => 
        \sample_filter_v2_out[6]\, sample_filter_v2_out_5 => 
        \sample_filter_v2_out[7]\, sample_filter_v2_out_6 => 
        \sample_filter_v2_out[8]\, sample_filter_v2_out_7 => 
        \sample_filter_v2_out[9]\, sample_filter_v2_out_8 => 
        \sample_filter_v2_out[10]\, sample_filter_v2_out_9 => 
        \sample_filter_v2_out[11]\, sample_filter_v2_out_10 => 
        \sample_filter_v2_out[12]\, sample_filter_v2_out_11 => 
        \sample_filter_v2_out[13]\, sample_filter_v2_out_12 => 
        \sample_filter_v2_out[14]\, sample_filter_v2_out_13 => 
        \sample_filter_v2_out[15]\, sample_filter_v2_out_14 => 
        \sample_filter_v2_out[16]\, sample_filter_v2_out_15 => 
        \sample_filter_v2_out[17]\, sample_filter_v2_out_18 => 
        \sample_filter_v2_out[20]\, sample_filter_v2_out_19 => 
        \sample_filter_v2_out[21]\, sample_filter_v2_out_20 => 
        \sample_filter_v2_out[22]\, sample_filter_v2_out_21 => 
        \sample_filter_v2_out[23]\, sample_filter_v2_out_22 => 
        \sample_filter_v2_out[24]\, sample_filter_v2_out_23 => 
        \sample_filter_v2_out[25]\, sample_filter_v2_out_24 => 
        \sample_filter_v2_out[26]\, sample_filter_v2_out_25 => 
        \sample_filter_v2_out[27]\, sample_filter_v2_out_26 => 
        \sample_filter_v2_out[28]\, sample_filter_v2_out_27 => 
        \sample_filter_v2_out[29]\, sample_filter_v2_out_28 => 
        \sample_filter_v2_out[30]\, sample_filter_v2_out_29 => 
        \sample_filter_v2_out[31]\, sample_filter_v2_out_30 => 
        \sample_filter_v2_out[32]\, sample_filter_v2_out_31 => 
        \sample_filter_v2_out[33]\, sample_filter_v2_out_32 => 
        \sample_filter_v2_out[34]\, sample_filter_v2_out_33 => 
        \sample_filter_v2_out[35]\, sample_filter_v2_out_36 => 
        \sample_filter_v2_out[38]\, sample_filter_v2_out_37 => 
        \sample_filter_v2_out[39]\, sample_filter_v2_out_38 => 
        \sample_filter_v2_out[40]\, sample_filter_v2_out_39 => 
        \sample_filter_v2_out[41]\, sample_filter_v2_out_40 => 
        \sample_filter_v2_out[42]\, sample_filter_v2_out_41 => 
        \sample_filter_v2_out[43]\, sample_filter_v2_out_42 => 
        \sample_filter_v2_out[44]\, sample_filter_v2_out_43 => 
        \sample_filter_v2_out[45]\, sample_filter_v2_out_44 => 
        \sample_filter_v2_out[46]\, sample_filter_v2_out_45 => 
        \sample_filter_v2_out[47]\, sample_filter_v2_out_46 => 
        \sample_filter_v2_out[48]\, sample_filter_v2_out_47 => 
        \sample_filter_v2_out[49]\, sample_filter_v2_out_48 => 
        \sample_filter_v2_out[50]\, sample_filter_v2_out_49 => 
        \sample_filter_v2_out[51]\, sample_filter_v2_out_50 => 
        \sample_filter_v2_out[52]\, sample_filter_v2_out_51 => 
        \sample_filter_v2_out[53]\, sample_filter_v2_out_54 => 
        \sample_filter_v2_out[56]\, sample_filter_v2_out_55 => 
        \sample_filter_v2_out[57]\, sample_filter_v2_out_56 => 
        \sample_filter_v2_out[58]\, sample_filter_v2_out_57 => 
        \sample_filter_v2_out[59]\, sample_filter_v2_out_58 => 
        \sample_filter_v2_out[60]\, sample_filter_v2_out_59 => 
        \sample_filter_v2_out[61]\, sample_filter_v2_out_60 => 
        \sample_filter_v2_out[62]\, sample_filter_v2_out_61 => 
        \sample_filter_v2_out[63]\, sample_filter_v2_out_62 => 
        \sample_filter_v2_out[64]\, sample_filter_v2_out_63 => 
        \sample_filter_v2_out[65]\, sample_filter_v2_out_64 => 
        \sample_filter_v2_out[66]\, sample_filter_v2_out_65 => 
        \sample_filter_v2_out[67]\, sample_filter_v2_out_66 => 
        \sample_filter_v2_out[68]\, sample_filter_v2_out_67 => 
        \sample_filter_v2_out[69]\, sample_filter_v2_out_68 => 
        \sample_filter_v2_out[70]\, sample_filter_v2_out_69 => 
        \sample_filter_v2_out[71]\, sample_filter_v2_out_90 => 
        \sample_filter_v2_out[92]\, sample_filter_v2_out_91 => 
        \sample_filter_v2_out[93]\, sample_filter_v2_out_92 => 
        \sample_filter_v2_out[94]\, sample_filter_v2_out_93 => 
        \sample_filter_v2_out[95]\, sample_filter_v2_out_94 => 
        \sample_filter_v2_out[96]\, sample_filter_v2_out_95 => 
        \sample_filter_v2_out[97]\, sample_filter_v2_out_96 => 
        \sample_filter_v2_out[98]\, sample_filter_v2_out_97 => 
        \sample_filter_v2_out[99]\, sample_filter_v2_out_98 => 
        \sample_filter_v2_out[100]\, sample_filter_v2_out_99 => 
        \sample_filter_v2_out[101]\, sample_filter_v2_out_100 => 
        \sample_filter_v2_out[102]\, sample_filter_v2_out_101 => 
        \sample_filter_v2_out[103]\, sample_filter_v2_out_102 => 
        \sample_filter_v2_out[104]\, sample_filter_v2_out_103 => 
        \sample_filter_v2_out[105]\, sample_filter_v2_out_104 => 
        \sample_filter_v2_out[106]\, sample_filter_v2_out_105 => 
        \sample_filter_v2_out[107]\, sample_filter_v2_out_108 => 
        \sample_filter_v2_out[110]\, sample_filter_v2_out_126 => 
        \sample_filter_v2_out[128]\, sample_filter_v2_out_109 => 
        \sample_filter_v2_out[111]\, sample_filter_v2_out_127 => 
        \sample_filter_v2_out[129]\, sample_filter_v2_out_110 => 
        \sample_filter_v2_out[112]\, sample_filter_v2_out_128 => 
        \sample_filter_v2_out[130]\, sample_filter_v2_out_111 => 
        \sample_filter_v2_out[113]\, sample_filter_v2_out_129 => 
        \sample_filter_v2_out[131]\, sample_filter_v2_out_112 => 
        \sample_filter_v2_out[114]\, sample_filter_v2_out_130 => 
        \sample_filter_v2_out[132]\, sample_filter_v2_out_113 => 
        \sample_filter_v2_out[115]\, sample_filter_v2_out_131 => 
        \sample_filter_v2_out[133]\, sample_filter_v2_out_114 => 
        \sample_filter_v2_out[116]\, sample_filter_v2_out_132 => 
        \sample_filter_v2_out[134]\, sample_filter_v2_out_115 => 
        \sample_filter_v2_out[117]\, sample_filter_v2_out_133 => 
        \sample_filter_v2_out[135]\, sample_filter_v2_out_116 => 
        \sample_filter_v2_out[118]\, sample_filter_v2_out_134 => 
        \sample_filter_v2_out[136]\, sample_filter_v2_out_117 => 
        \sample_filter_v2_out[119]\, sample_filter_v2_out_135 => 
        \sample_filter_v2_out[137]\, sample_filter_v2_out_118 => 
        \sample_filter_v2_out[120]\, sample_filter_v2_out_136 => 
        \sample_filter_v2_out[138]\, sample_filter_v2_out_119 => 
        \sample_filter_v2_out[121]\, sample_filter_v2_out_137 => 
        \sample_filter_v2_out[139]\, sample_filter_v2_out_120 => 
        \sample_filter_v2_out[122]\, sample_filter_v2_out_138 => 
        \sample_filter_v2_out[140]\, sample_filter_v2_out_121 => 
        \sample_filter_v2_out[123]\, sample_filter_v2_out_139 => 
        \sample_filter_v2_out[141]\, sample_filter_v2_out_122 => 
        \sample_filter_v2_out[124]\, sample_filter_v2_out_140 => 
        \sample_filter_v2_out[142]\, sample_filter_v2_out_123 => 
        \sample_filter_v2_out[125]\, sample_filter_v2_out_141 => 
        \sample_filter_v2_out[143]\, sample_6(15) => 
        \sample_6[15]\, sample_6(14) => \sample_6[14]\, 
        sample_6(13) => \sample_6[13]\, sample_6(12) => 
        \sample_6[12]\, sample_6(11) => \sample_6[11]\, 
        sample_6(10) => \sample_6[10]\, sample_6(9) => 
        \sample_6[9]\, sample_6(8) => \sample_6[8]\, sample_6(7)
         => \sample_6[7]\, sample_6(6) => \sample_6[6]\, 
        sample_6(5) => \sample_6[5]\, sample_6(4) => 
        \sample_6[4]\, sample_6(3) => \sample_6[3]\, sample_6(2)
         => \sample_6[2]\, sample_6(1) => \sample_6[1]\, 
        sample_6(0) => \sample_6[0]\, sample_5(15) => 
        \sample_5[15]\, sample_5(14) => \sample_5[14]\, 
        sample_5(13) => \sample_5[13]\, sample_5(12) => 
        \sample_5[12]\, sample_5(11) => \sample_5[11]\, 
        sample_5(10) => \sample_5[10]\, sample_5(9) => 
        \sample_5[9]\, sample_5(8) => \sample_5[8]\, sample_5(7)
         => \sample_5[7]\, sample_5(6) => \sample_5[6]\, 
        sample_5(5) => \sample_5[5]\, sample_5(4) => 
        \sample_5[4]\, sample_5(3) => \sample_5[3]\, sample_5(2)
         => \sample_5[2]\, sample_5(1) => \sample_5[1]\, 
        sample_5(0) => \sample_5[0]\, sample_2(15) => 
        \sample_2[15]\, sample_2(14) => \sample_2[14]\, 
        sample_2(13) => \sample_2[13]\, sample_2(12) => 
        \sample_2[12]\, sample_2(11) => \sample_2[11]\, 
        sample_2(10) => \sample_2[10]\, sample_2(9) => 
        \sample_2[9]\, sample_2(8) => \sample_2[8]\, sample_2(7)
         => \sample_2[7]\, sample_2(6) => \sample_2[6]\, 
        sample_2(5) => \sample_2[5]\, sample_2(4) => 
        \sample_2[4]\, sample_2(3) => \sample_2[3]\, sample_2(2)
         => \sample_2[2]\, sample_2(1) => \sample_2[1]\, 
        sample_2(0) => \sample_2[0]\, sample_0(15) => 
        \sample_0[15]\, sample_0(14) => \sample_0[14]\, 
        sample_0(13) => \sample_0[13]\, sample_0(12) => 
        \sample_0[12]\, sample_0(11) => \sample_0[11]\, 
        sample_0(10) => \sample_0[10]\, sample_0(9) => 
        \sample_0[9]\, sample_0(8) => \sample_0[8]\, sample_0(7)
         => \sample_0[7]\, sample_0(6) => \sample_0[6]\, 
        sample_0(5) => \sample_0[5]\, sample_0(4) => 
        \sample_0[4]\, sample_0(3) => \sample_0[3]\, sample_0(2)
         => \sample_0[2]\, sample_0(1) => \sample_0[1]\, 
        sample_0(0) => \sample_0[0]\, sample_1(15) => 
        \sample_1[15]\, sample_1(14) => \sample_1[14]\, 
        sample_1(13) => \sample_1[13]\, sample_1(12) => 
        \sample_1[12]\, sample_1(11) => \sample_1[11]\, 
        sample_1(10) => \sample_1[10]\, sample_1(9) => 
        \sample_1[9]\, sample_1(8) => \sample_1[8]\, sample_1(7)
         => \sample_1[7]\, sample_1(6) => \sample_1[6]\, 
        sample_1(5) => \sample_1[5]\, sample_1(4) => 
        \sample_1[4]\, sample_1(3) => \sample_1[3]\, sample_1(2)
         => \sample_1[2]\, sample_1(1) => \sample_1[1]\, 
        sample_1(0) => \sample_1[0]\, sample_3(15) => 
        \sample_3[15]\, sample_3(14) => \sample_3[14]\, 
        sample_3(13) => \sample_3[13]\, sample_3(12) => 
        \sample_3[12]\, sample_3(11) => \sample_3[11]\, 
        sample_3(10) => \sample_3[10]\, sample_3(9) => 
        \sample_3[9]\, sample_3(8) => \sample_3[8]\, sample_3(7)
         => \sample_3[7]\, sample_3(6) => \sample_3[6]\, 
        sample_3(5) => \sample_3[5]\, sample_3(4) => 
        \sample_3[4]\, sample_3(3) => \sample_3[3]\, sample_3(2)
         => \sample_3[2]\, sample_3(1) => \sample_3[1]\, 
        sample_3(0) => \sample_3[0]\, sample_4(15) => 
        \sample_4[15]\, sample_4(14) => \sample_4[14]\, 
        sample_4(13) => \sample_4[13]\, sample_4(12) => 
        \sample_4[12]\, sample_4(11) => \sample_4[11]\, 
        sample_4(10) => \sample_4[10]\, sample_4(9) => 
        \sample_4[9]\, sample_4(8) => \sample_4[8]\, sample_4(7)
         => \sample_4[7]\, sample_4(6) => \sample_4[6]\, 
        sample_4(5) => \sample_4[5]\, sample_4(4) => 
        \sample_4[4]\, sample_4(3) => \sample_4[3]\, sample_4(2)
         => \sample_4[2]\, sample_4(1) => \sample_4[1]\, 
        sample_4(0) => \sample_4[0]\, sample_7(15) => 
        \sample_7[15]\, sample_7(14) => \sample_7[14]\, 
        sample_7(13) => \sample_7[13]\, sample_7(12) => 
        \sample_7[12]\, sample_7(11) => \sample_7[11]\, 
        sample_7(10) => \sample_7[10]\, sample_7(9) => 
        \sample_7[9]\, sample_7(8) => \sample_7[8]\, sample_7(7)
         => \sample_7[7]\, sample_7(6) => \sample_7[6]\, 
        sample_7(5) => \sample_7[5]\, sample_7(4) => 
        \sample_7[4]\, sample_7(3) => \sample_7[3]\, sample_7(2)
         => \sample_7[2]\, sample_7(1) => \sample_7[1]\, 
        sample_7(0) => \sample_7[0]\, IIR_CEL_CTRLR_v2_VCC => 
        lpp_top_lfr_wf_picker_ip_VCC, IIR_CEL_CTRLR_v2_GND => 
        lpp_top_lfr_wf_picker_ip_GND, HRESETn_c => HRESETn_c, 
        HCLK_c => HCLK_c, sample_filter_v2_out_val => 
        sample_filter_v2_out_val, sample_val_delay => 
        \sample_val_delay\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I101_Y_0 : 
        XNOR2
      port map(A => N288_i, B => N195, Y => 
        \sample_data_shaping_f1_f0_s[8]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[103]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_113[103]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[103]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I22_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[137]\, B => 
        \sample_filter_v2_out[119]\, Y => N191);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[135]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[135]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[135]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I98_Y_0 : 
        AX1D
      port map(A => I85_un1_Y, B => N274_0, C => N189, Y => 
        \sample_data_shaping_f1_f0_s[5]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I24_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[135]\, B => 
        \sample_filter_v2_out[117]\, Y => N195);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[28]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[28]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[28]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out_RNO[110]\ : 
        MX2
      port map(A => \sample_filter_v2_out[110]\, B => 
        \sample_data_shaping_f1_f0_s[15]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_373[110]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I108_Y_0 : 
        XNOR3
      port map(A => \sample_filter_v2_out[110]\, B => 
        \sample_filter_v2_out[128]\, C => N240, Y => 
        \sample_data_shaping_f1_f0_s[15]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I78_Y : 
        AO1
      port map(A => N268, B => N265, C => N264, Y => N270);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I71_Y : 
        AO1C
      port map(A => N255, B => N258, C => N254_0, Y => N260);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I49_Y_0 : 
        AO18
      port map(A => N198_0, B => \sample_filter_v2_out[133]\, C
         => \sample_filter_v2_out[115]\, Y => 
        SUB_16x16_medium_area_I49_Y_0_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I17_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[124]\, B => 
        \sample_filter_v2_out[106]\, Y => N181_0);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[30]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[30]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[30]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I33_Y : 
        XAI1A
      port map(A => \sample_filter_v2_out[111]\, B => 
        \sample_filter_v2_out[129]\, C => N205, Y => N212_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I17_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[124]\, B => 
        \sample_filter_v2_out[142]\, Y => N182_0);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I104_Y_0 : 
        XOR2
      port map(A => N258, B => N201, Y => 
        \sample_data_shaping_f1_f0_s[11]\);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[119]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_157[119]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[119]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I49_Y_0 : 
        AO18
      port map(A => N198, B => \sample_filter_v2_out[115]\, C => 
        \sample_filter_v2_out[97]\, Y => 
        SUB_16x16_medium_area_I49_Y_0);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out_RNO[101]\ : 
        MX2
      port map(A => \sample_filter_v2_out[101]\, B => 
        \sample_data_shaping_f2_f1_s[6]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_161[101]\);
    
    sample_val_delay_RNI8T43 : CLKINT
      port map(A => sample_val_delay_0, Y => \sample_val_delay\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I29_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[94]\, B => 
        \sample_filter_v2_out[112]\, Y => N206);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out_RNO[93]\ : 
        MX2
      port map(A => \sample_filter_v2_out[93]\, B => 
        \sample_data_shaping_f2_f1_s[14]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_353[93]\);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[47]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[47]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[47]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[120]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_133[120]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[120]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[13]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[13]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[13]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[32]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[32]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[32]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I21_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[102]\, B => 
        \sample_filter_v2_out[120]\, Y => N190);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[15]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[15]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[15]\);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out_RNO[95]\ : 
        MX2
      port map(A => \sample_filter_v2_out[95]\, B => 
        \sample_data_shaping_f2_f1_s[12]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_305[95]\);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[113]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_301[113]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[113]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I56_Y_1 : 
        AOI1B
      port map(A => N274_0, B => N220_0, C => 
        SUB_16x16_medium_area_I56_Y_0_0, Y => 
        SUB_16x16_medium_area_I56_Y_1_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I20_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[121]\, B => 
        \sample_filter_v2_out[103]\, Y => N187_0);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out_RNO[123]\ : 
        MX2
      port map(A => \sample_filter_v2_out[123]\, B => 
        \sample_data_shaping_f1_f0_s[2]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_61[123]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[67]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[67]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[67]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I87_un1_Y : 
        OA1A
      port map(A => I64_un1_Y, B => N244, C => N201_0, Y => 
        SUB_16x16_medium_area_I87_un1_Y);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I71_un1_Y : 
        OA1A
      port map(A => I64_un1_Y, B => N244, C => N255_0, Y => 
        I71_un1_Y);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I37_Y : 
        NOR2B
      port map(A => N199, B => N197_0, Y => N216_0);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[104]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_89[104]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[104]\);
    
    sample_val_delay : DFN1C0
      port map(D => sample_val, CLK => HCLK_c, CLR => HRESETn_c, 
        Q => sample_val_delay_0);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[35]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[35]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[35]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I48_Y : 
        NOR2B
      port map(A => N255_0, B => N212, Y => N229);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I57_un1_Y_0 : 
        NOR2B
      port map(A => N229, B => N245, Y => 
        SUB_16x16_medium_area_I57_un1_Y_0);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[129]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[129]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[129]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I94_Y_0 : 
        XOR2
      port map(A => N225_0, B => N181, Y => 
        \sample_data_shaping_f1_f0_s[1]\);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[107]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_17[107]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[107]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I28_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[113]\, B => 
        \sample_filter_v2_out[95]\, Y => N203);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I107_Y_0 : 
        XNOR3
      port map(A => \sample_filter_v2_out[111]\, B => 
        \sample_filter_v2_out[129]\, C => N282_i, Y => 
        \sample_data_shaping_f1_f0_s_i[14]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I19_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[140]\, B => 
        \sample_filter_v2_out[122]\, Y => N185);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[137]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[137]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[137]\);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[11]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[11]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[11]\);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[46]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[46]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[46]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[110]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_373[110]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[110]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[61]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[61]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[61]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I102_Y_0 : 
        XOR2
      port map(A => N270, B => N197, Y => 
        \sample_data_shaping_f1_f0_s[9]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[68]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[68]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[68]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I42_Y : 
        AO13
      port map(A => N186_0, B => \sample_filter_v2_out[103]\, C
         => \sample_filter_v2_out[121]\, Y => N274);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[57]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[57]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[57]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I107_Y_0 : 
        AX1D
      port map(A => I86_un1_Y, B => N206, C => N207, Y => 
        \sample_data_shaping_f2_f1_s[14]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I53_un1_Y_0 : 
        XA1A
      port map(A => \sample_filter_v2_out[105]\, B => 
        \sample_filter_v2_out[123]\, C => N225, Y => 
        SUB_16x16_medium_area_I53_un1_Y_0);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[49]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[49]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[49]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out_RNO[104]\ : 
        MX2
      port map(A => \sample_filter_v2_out[104]\, B => 
        \sample_data_shaping_f2_f1_s[3]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_89[104]\);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[17]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[17]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[17]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I92_Y : 
        AO18
      port map(A => N225, B => \sample_filter_v2_out[124]\, C => 
        \sample_filter_v2_out[106]\, Y => N294_i);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I105_Y_0 : 
        XOR3
      port map(A => \sample_filter_v2_out[113]\, B => 
        \sample_filter_v2_out[131]\, C => N284_i, Y => 
        \sample_data_shaping_f1_f0_s[12]\);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out_RNO[116]\ : 
        MX2
      port map(A => \sample_filter_v2_out[116]\, B => 
        \sample_data_shaping_f1_f0_s[9]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_229[116]\);
    
    Downsampling_f3 : Downsampling_6_16_256
      port map(sample_f1(111) => \sample_f1[111]\, sample_f1(110)
         => \sample_f1[110]\, sample_f1(109) => \sample_f1[109]\, 
        sample_f1(108) => \sample_f1[108]\, sample_f1(107) => 
        \sample_f1[107]\, sample_f1(106) => \sample_f1[106]\, 
        sample_f1(105) => \sample_f1[105]\, sample_f1(104) => 
        \sample_f1[104]\, sample_f1(103) => \sample_f1[103]\, 
        sample_f1(102) => \sample_f1[102]\, sample_f1(101) => 
        \sample_f1[101]\, sample_f1(100) => \sample_f1[100]\, 
        sample_f1(99) => \sample_f1[99]\, sample_f1(98) => 
        \sample_f1[98]\, sample_f1(97) => \sample_f1[97]\, 
        sample_f1(96) => \sample_f1[96]\, sample_f1(95) => 
        \sample_f1[95]\, sample_f1(94) => \sample_f1[94]\, 
        sample_f1(93) => \sample_f1[93]\, sample_f1(92) => 
        \sample_f1[92]\, sample_f1(91) => \sample_f1[91]\, 
        sample_f1(90) => \sample_f1[90]\, sample_f1(89) => 
        \sample_f1[89]\, sample_f1(88) => \sample_f1[88]\, 
        sample_f1(87) => \sample_f1[87]\, sample_f1(86) => 
        \sample_f1[86]\, sample_f1(85) => \sample_f1[85]\, 
        sample_f1(84) => \sample_f1[84]\, sample_f1(83) => 
        \sample_f1[83]\, sample_f1(82) => \sample_f1[82]\, 
        sample_f1(81) => \sample_f1[81]\, sample_f1(80) => 
        \sample_f1[80]\, sample_f1_wdata_95 => 
        \sample_f1_wdata[95]\, sample_f1_wdata_94 => 
        \sample_f1_wdata[94]\, sample_f1_wdata_93 => 
        \sample_f1_wdata[93]\, sample_f1_wdata_92 => 
        \sample_f1_wdata[92]\, sample_f1_wdata_91 => 
        \sample_f1_wdata[91]\, sample_f1_wdata_90 => 
        \sample_f1_wdata[90]\, sample_f1_wdata_89 => 
        \sample_f1_wdata[89]\, sample_f1_wdata_88 => 
        \sample_f1_wdata[88]\, sample_f1_wdata_87 => 
        \sample_f1_wdata[87]\, sample_f1_wdata_86 => 
        \sample_f1_wdata[86]\, sample_f1_wdata_85 => 
        \sample_f1_wdata[85]\, sample_f1_wdata_84 => 
        \sample_f1_wdata[84]\, sample_f1_wdata_83 => 
        \sample_f1_wdata[83]\, sample_f1_wdata_82 => 
        \sample_f1_wdata[82]\, sample_f1_wdata_81 => 
        \sample_f1_wdata[81]\, sample_f1_wdata_80 => 
        \sample_f1_wdata[80]\, sample_f1_wdata_79 => 
        \sample_f1_wdata[79]\, sample_f1_wdata_78 => 
        \sample_f1_wdata[78]\, sample_f1_wdata_77 => 
        \sample_f1_wdata[77]\, sample_f1_wdata_76 => 
        \sample_f1_wdata[76]\, sample_f1_wdata_75 => 
        \sample_f1_wdata[75]\, sample_f1_wdata_74 => 
        \sample_f1_wdata[74]\, sample_f1_wdata_73 => 
        \sample_f1_wdata[73]\, sample_f1_wdata_72 => 
        \sample_f1_wdata[72]\, sample_f1_wdata_71 => 
        \sample_f1_wdata[71]\, sample_f1_wdata_70 => 
        \sample_f1_wdata[70]\, sample_f1_wdata_69 => 
        \sample_f1_wdata[69]\, sample_f1_wdata_68 => 
        \sample_f1_wdata[68]\, sample_f1_wdata_67 => 
        \sample_f1_wdata[67]\, sample_f1_wdata_66 => 
        \sample_f1_wdata[66]\, sample_f1_wdata_65 => 
        \sample_f1_wdata[65]\, sample_f1_wdata_64 => 
        \sample_f1_wdata[64]\, sample_f1_wdata_63 => 
        \sample_f1_wdata[63]\, sample_f1_wdata_62 => 
        \sample_f1_wdata[62]\, sample_f1_wdata_61 => 
        \sample_f1_wdata[61]\, sample_f1_wdata_60 => 
        \sample_f1_wdata[60]\, sample_f1_wdata_59 => 
        \sample_f1_wdata[59]\, sample_f1_wdata_58 => 
        \sample_f1_wdata[58]\, sample_f1_wdata_57 => 
        \sample_f1_wdata[57]\, sample_f1_wdata_56 => 
        \sample_f1_wdata[56]\, sample_f1_wdata_55 => 
        \sample_f1_wdata[55]\, sample_f1_wdata_54 => 
        \sample_f1_wdata[54]\, sample_f1_wdata_53 => 
        \sample_f1_wdata[53]\, sample_f1_wdata_52 => 
        \sample_f1_wdata[52]\, sample_f1_wdata_51 => 
        \sample_f1_wdata[51]\, sample_f1_wdata_50 => 
        \sample_f1_wdata[50]\, sample_f1_wdata_49 => 
        \sample_f1_wdata[49]\, sample_f1_wdata_48 => 
        \sample_f1_wdata[48]\, sample_f1_wdata_15 => 
        \sample_f1_wdata[15]\, sample_f1_wdata_14 => 
        \sample_f1_wdata[14]\, sample_f1_wdata_13 => 
        \sample_f1_wdata[13]\, sample_f1_wdata_12 => 
        \sample_f1_wdata[12]\, sample_f1_wdata_11 => 
        \sample_f1_wdata[11]\, sample_f1_wdata_10 => 
        \sample_f1_wdata[10]\, sample_f1_wdata_9 => 
        \sample_f1_wdata[9]\, sample_f1_wdata_8 => 
        \sample_f1_wdata[8]\, sample_f1_wdata_7 => 
        \sample_f1_wdata[7]\, sample_f1_wdata_6 => 
        \sample_f1_wdata[6]\, sample_f1_wdata_5 => 
        \sample_f1_wdata[5]\, sample_f1_wdata_4 => 
        \sample_f1_wdata[4]\, sample_f1_wdata_3 => 
        \sample_f1_wdata[3]\, sample_f1_wdata_2 => 
        \sample_f1_wdata[2]\, sample_f1_wdata_1 => 
        \sample_f1_wdata[1]\, sample_f1_wdata_0 => 
        \sample_f1_wdata[0]\, sample_f3_wdata(95) => 
        \sample_f3_wdata[95]\, sample_f3_wdata(94) => 
        \sample_f3_wdata[94]\, sample_f3_wdata(93) => 
        \sample_f3_wdata[93]\, sample_f3_wdata(92) => 
        \sample_f3_wdata[92]\, sample_f3_wdata(91) => 
        \sample_f3_wdata[91]\, sample_f3_wdata(90) => 
        \sample_f3_wdata[90]\, sample_f3_wdata(89) => 
        \sample_f3_wdata[89]\, sample_f3_wdata(88) => 
        \sample_f3_wdata[88]\, sample_f3_wdata(87) => 
        \sample_f3_wdata[87]\, sample_f3_wdata(86) => 
        \sample_f3_wdata[86]\, sample_f3_wdata(85) => 
        \sample_f3_wdata[85]\, sample_f3_wdata(84) => 
        \sample_f3_wdata[84]\, sample_f3_wdata(83) => 
        \sample_f3_wdata[83]\, sample_f3_wdata(82) => 
        \sample_f3_wdata[82]\, sample_f3_wdata(81) => 
        \sample_f3_wdata[81]\, sample_f3_wdata(80) => 
        \sample_f3_wdata[80]\, sample_f3_wdata(79) => 
        \sample_f3_wdata[79]\, sample_f3_wdata(78) => 
        \sample_f3_wdata[78]\, sample_f3_wdata(77) => 
        \sample_f3_wdata[77]\, sample_f3_wdata(76) => 
        \sample_f3_wdata[76]\, sample_f3_wdata(75) => 
        \sample_f3_wdata[75]\, sample_f3_wdata(74) => 
        \sample_f3_wdata[74]\, sample_f3_wdata(73) => 
        \sample_f3_wdata[73]\, sample_f3_wdata(72) => 
        \sample_f3_wdata[72]\, sample_f3_wdata(71) => 
        \sample_f3_wdata[71]\, sample_f3_wdata(70) => 
        \sample_f3_wdata[70]\, sample_f3_wdata(69) => 
        \sample_f3_wdata[69]\, sample_f3_wdata(68) => 
        \sample_f3_wdata[68]\, sample_f3_wdata(67) => 
        \sample_f3_wdata[67]\, sample_f3_wdata(66) => 
        \sample_f3_wdata[66]\, sample_f3_wdata(65) => 
        \sample_f3_wdata[65]\, sample_f3_wdata(64) => 
        \sample_f3_wdata[64]\, sample_f3_wdata(63) => 
        \sample_f3_wdata[63]\, sample_f3_wdata(62) => 
        \sample_f3_wdata[62]\, sample_f3_wdata(61) => 
        \sample_f3_wdata[61]\, sample_f3_wdata(60) => 
        \sample_f3_wdata[60]\, sample_f3_wdata(59) => 
        \sample_f3_wdata[59]\, sample_f3_wdata(58) => 
        \sample_f3_wdata[58]\, sample_f3_wdata(57) => 
        \sample_f3_wdata[57]\, sample_f3_wdata(56) => 
        \sample_f3_wdata[56]\, sample_f3_wdata(55) => 
        \sample_f3_wdata[55]\, sample_f3_wdata(54) => 
        \sample_f3_wdata[54]\, sample_f3_wdata(53) => 
        \sample_f3_wdata[53]\, sample_f3_wdata(52) => 
        \sample_f3_wdata[52]\, sample_f3_wdata(51) => 
        \sample_f3_wdata[51]\, sample_f3_wdata(50) => 
        \sample_f3_wdata[50]\, sample_f3_wdata(49) => 
        \sample_f3_wdata[49]\, sample_f3_wdata(48) => 
        \sample_f3_wdata[48]\, sample_f3_wdata(47) => 
        \sample_f3_wdata[47]\, sample_f3_wdata(46) => 
        \sample_f3_wdata[46]\, sample_f3_wdata(45) => 
        \sample_f3_wdata[45]\, sample_f3_wdata(44) => 
        \sample_f3_wdata[44]\, sample_f3_wdata(43) => 
        \sample_f3_wdata[43]\, sample_f3_wdata(42) => 
        \sample_f3_wdata[42]\, sample_f3_wdata(41) => 
        \sample_f3_wdata[41]\, sample_f3_wdata(40) => 
        \sample_f3_wdata[40]\, sample_f3_wdata(39) => 
        \sample_f3_wdata[39]\, sample_f3_wdata(38) => 
        \sample_f3_wdata[38]\, sample_f3_wdata(37) => 
        \sample_f3_wdata[37]\, sample_f3_wdata(36) => 
        \sample_f3_wdata[36]\, sample_f3_wdata(35) => 
        \sample_f3_wdata[35]\, sample_f3_wdata(34) => 
        \sample_f3_wdata[34]\, sample_f3_wdata(33) => 
        \sample_f3_wdata[33]\, sample_f3_wdata(32) => 
        \sample_f3_wdata[32]\, sample_f3_wdata(31) => 
        \sample_f3_wdata[31]\, sample_f3_wdata(30) => 
        \sample_f3_wdata[30]\, sample_f3_wdata(29) => 
        \sample_f3_wdata[29]\, sample_f3_wdata(28) => 
        \sample_f3_wdata[28]\, sample_f3_wdata(27) => 
        \sample_f3_wdata[27]\, sample_f3_wdata(26) => 
        \sample_f3_wdata[26]\, sample_f3_wdata(25) => 
        \sample_f3_wdata[25]\, sample_f3_wdata(24) => 
        \sample_f3_wdata[24]\, sample_f3_wdata(23) => 
        \sample_f3_wdata[23]\, sample_f3_wdata(22) => 
        \sample_f3_wdata[22]\, sample_f3_wdata(21) => 
        \sample_f3_wdata[21]\, sample_f3_wdata(20) => 
        \sample_f3_wdata[20]\, sample_f3_wdata(19) => 
        \sample_f3_wdata[19]\, sample_f3_wdata(18) => 
        \sample_f3_wdata[18]\, sample_f3_wdata(17) => 
        \sample_f3_wdata[17]\, sample_f3_wdata(16) => 
        \sample_f3_wdata[16]\, sample_f3_wdata(15) => 
        \sample_f3_wdata[15]\, sample_f3_wdata(14) => 
        \sample_f3_wdata[14]\, sample_f3_wdata(13) => 
        \sample_f3_wdata[13]\, sample_f3_wdata(12) => 
        \sample_f3_wdata[12]\, sample_f3_wdata(11) => 
        \sample_f3_wdata[11]\, sample_f3_wdata(10) => 
        \sample_f3_wdata[10]\, sample_f3_wdata(9) => 
        \sample_f3_wdata[9]\, sample_f3_wdata(8) => 
        \sample_f3_wdata[8]\, sample_f3_wdata(7) => 
        \sample_f3_wdata[7]\, sample_f3_wdata(6) => 
        \sample_f3_wdata[6]\, sample_f3_wdata(5) => 
        \sample_f3_wdata[5]\, sample_f3_wdata(4) => 
        \sample_f3_wdata[4]\, sample_f3_wdata(3) => 
        \sample_f3_wdata[3]\, sample_f3_wdata(2) => 
        \sample_f3_wdata[2]\, sample_f3_wdata(1) => 
        \sample_f3_wdata[1]\, sample_f3_wdata(0) => 
        \sample_f3_wdata[0]\, sample_f1_val => sample_f1_val, 
        HCLK_c => HCLK_c, sample_f3_val => sample_f3_val, 
        HRESETn_c => HRESETn_c, sample_f1_val_0 => 
        sample_f1_val_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I34_Y : 
        AO18
      port map(A => N202, B => \sample_filter_v2_out[131]\, C => 
        \sample_filter_v2_out[113]\, Y => N254_0);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out_RNO[115]\ : 
        MX2
      port map(A => \sample_filter_v2_out[115]\, B => 
        \sample_data_shaping_f1_f0_s[10]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_253[115]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    Downsampling_f2 : Downsampling_6_16_96
      port map(sample_f0(111) => \sample_f0[111]\, sample_f0(110)
         => \sample_f0[110]\, sample_f0(109) => \sample_f0[109]\, 
        sample_f0(108) => \sample_f0[108]\, sample_f0(107) => 
        \sample_f0[107]\, sample_f0(106) => \sample_f0[106]\, 
        sample_f0(105) => \sample_f0[105]\, sample_f0(104) => 
        \sample_f0[104]\, sample_f0(103) => \sample_f0[103]\, 
        sample_f0(102) => \sample_f0[102]\, sample_f0(101) => 
        \sample_f0[101]\, sample_f0(100) => \sample_f0[100]\, 
        sample_f0(99) => \sample_f0[99]\, sample_f0(98) => 
        \sample_f0[98]\, sample_f0(97) => \sample_f0[97]\, 
        sample_f0(96) => \sample_f0[96]\, sample_f0(95) => 
        \sample_f0[95]\, sample_f0(94) => \sample_f0[94]\, 
        sample_f0(93) => \sample_f0[93]\, sample_f0(92) => 
        \sample_f0[92]\, sample_f0(91) => \sample_f0[91]\, 
        sample_f0(90) => \sample_f0[90]\, sample_f0(89) => 
        \sample_f0[89]\, sample_f0(88) => \sample_f0[88]\, 
        sample_f0(87) => \sample_f0[87]\, sample_f0(86) => 
        \sample_f0[86]\, sample_f0(85) => \sample_f0[85]\, 
        sample_f0(84) => \sample_f0[84]\, sample_f0(83) => 
        \sample_f0[83]\, sample_f0(82) => \sample_f0[82]\, 
        sample_f0(81) => \sample_f0[81]\, sample_f0(80) => 
        \sample_f0[80]\, sample_f0_wdata_95 => 
        \sample_f0_wdata[95]\, sample_f0_wdata_94 => 
        \sample_f0_wdata[94]\, sample_f0_wdata_93 => 
        \sample_f0_wdata[93]\, sample_f0_wdata_92 => 
        \sample_f0_wdata[92]\, sample_f0_wdata_91 => 
        \sample_f0_wdata[91]\, sample_f0_wdata_90 => 
        \sample_f0_wdata[90]\, sample_f0_wdata_89 => 
        \sample_f0_wdata[89]\, sample_f0_wdata_88 => 
        \sample_f0_wdata[88]\, sample_f0_wdata_87 => 
        \sample_f0_wdata[87]\, sample_f0_wdata_86 => 
        \sample_f0_wdata[86]\, sample_f0_wdata_85 => 
        \sample_f0_wdata[85]\, sample_f0_wdata_84 => 
        \sample_f0_wdata[84]\, sample_f0_wdata_83 => 
        \sample_f0_wdata[83]\, sample_f0_wdata_82 => 
        \sample_f0_wdata[82]\, sample_f0_wdata_81 => 
        \sample_f0_wdata[81]\, sample_f0_wdata_80 => 
        \sample_f0_wdata[80]\, sample_f0_wdata_79 => 
        \sample_f0_wdata[79]\, sample_f0_wdata_78 => 
        \sample_f0_wdata[78]\, sample_f0_wdata_77 => 
        \sample_f0_wdata[77]\, sample_f0_wdata_76 => 
        \sample_f0_wdata[76]\, sample_f0_wdata_75 => 
        \sample_f0_wdata[75]\, sample_f0_wdata_74 => 
        \sample_f0_wdata[74]\, sample_f0_wdata_73 => 
        \sample_f0_wdata[73]\, sample_f0_wdata_72 => 
        \sample_f0_wdata[72]\, sample_f0_wdata_71 => 
        \sample_f0_wdata[71]\, sample_f0_wdata_70 => 
        \sample_f0_wdata[70]\, sample_f0_wdata_69 => 
        \sample_f0_wdata[69]\, sample_f0_wdata_68 => 
        \sample_f0_wdata[68]\, sample_f0_wdata_67 => 
        \sample_f0_wdata[67]\, sample_f0_wdata_66 => 
        \sample_f0_wdata[66]\, sample_f0_wdata_65 => 
        \sample_f0_wdata[65]\, sample_f0_wdata_64 => 
        \sample_f0_wdata[64]\, sample_f0_wdata_63 => 
        \sample_f0_wdata[63]\, sample_f0_wdata_62 => 
        \sample_f0_wdata[62]\, sample_f0_wdata_61 => 
        \sample_f0_wdata[61]\, sample_f0_wdata_60 => 
        \sample_f0_wdata[60]\, sample_f0_wdata_59 => 
        \sample_f0_wdata[59]\, sample_f0_wdata_58 => 
        \sample_f0_wdata[58]\, sample_f0_wdata_57 => 
        \sample_f0_wdata[57]\, sample_f0_wdata_56 => 
        \sample_f0_wdata[56]\, sample_f0_wdata_55 => 
        \sample_f0_wdata[55]\, sample_f0_wdata_54 => 
        \sample_f0_wdata[54]\, sample_f0_wdata_53 => 
        \sample_f0_wdata[53]\, sample_f0_wdata_52 => 
        \sample_f0_wdata[52]\, sample_f0_wdata_51 => 
        \sample_f0_wdata[51]\, sample_f0_wdata_50 => 
        \sample_f0_wdata[50]\, sample_f0_wdata_49 => 
        \sample_f0_wdata[49]\, sample_f0_wdata_48 => 
        \sample_f0_wdata[48]\, sample_f0_wdata_15 => 
        \sample_f0_wdata[15]\, sample_f0_wdata_14 => 
        \sample_f0_wdata[14]\, sample_f0_wdata_13 => 
        \sample_f0_wdata[13]\, sample_f0_wdata_12 => 
        \sample_f0_wdata[12]\, sample_f0_wdata_11 => 
        \sample_f0_wdata[11]\, sample_f0_wdata_10 => 
        \sample_f0_wdata[10]\, sample_f0_wdata_9 => 
        \sample_f0_wdata[9]\, sample_f0_wdata_8 => 
        \sample_f0_wdata[8]\, sample_f0_wdata_7 => 
        \sample_f0_wdata[7]\, sample_f0_wdata_6 => 
        \sample_f0_wdata[6]\, sample_f0_wdata_5 => 
        \sample_f0_wdata[5]\, sample_f0_wdata_4 => 
        \sample_f0_wdata[4]\, sample_f0_wdata_3 => 
        \sample_f0_wdata[3]\, sample_f0_wdata_2 => 
        \sample_f0_wdata[2]\, sample_f0_wdata_1 => 
        \sample_f0_wdata[1]\, sample_f0_wdata_0 => 
        \sample_f0_wdata[0]\, sample_f2_wdata(95) => 
        \sample_f2_wdata[95]\, sample_f2_wdata(94) => 
        \sample_f2_wdata[94]\, sample_f2_wdata(93) => 
        \sample_f2_wdata[93]\, sample_f2_wdata(92) => 
        \sample_f2_wdata[92]\, sample_f2_wdata(91) => 
        \sample_f2_wdata[91]\, sample_f2_wdata(90) => 
        \sample_f2_wdata[90]\, sample_f2_wdata(89) => 
        \sample_f2_wdata[89]\, sample_f2_wdata(88) => 
        \sample_f2_wdata[88]\, sample_f2_wdata(87) => 
        \sample_f2_wdata[87]\, sample_f2_wdata(86) => 
        \sample_f2_wdata[86]\, sample_f2_wdata(85) => 
        \sample_f2_wdata[85]\, sample_f2_wdata(84) => 
        \sample_f2_wdata[84]\, sample_f2_wdata(83) => 
        \sample_f2_wdata[83]\, sample_f2_wdata(82) => 
        \sample_f2_wdata[82]\, sample_f2_wdata(81) => 
        \sample_f2_wdata[81]\, sample_f2_wdata(80) => 
        \sample_f2_wdata[80]\, sample_f2_wdata(79) => 
        \sample_f2_wdata[79]\, sample_f2_wdata(78) => 
        \sample_f2_wdata[78]\, sample_f2_wdata(77) => 
        \sample_f2_wdata[77]\, sample_f2_wdata(76) => 
        \sample_f2_wdata[76]\, sample_f2_wdata(75) => 
        \sample_f2_wdata[75]\, sample_f2_wdata(74) => 
        \sample_f2_wdata[74]\, sample_f2_wdata(73) => 
        \sample_f2_wdata[73]\, sample_f2_wdata(72) => 
        \sample_f2_wdata[72]\, sample_f2_wdata(71) => 
        \sample_f2_wdata[71]\, sample_f2_wdata(70) => 
        \sample_f2_wdata[70]\, sample_f2_wdata(69) => 
        \sample_f2_wdata[69]\, sample_f2_wdata(68) => 
        \sample_f2_wdata[68]\, sample_f2_wdata(67) => 
        \sample_f2_wdata[67]\, sample_f2_wdata(66) => 
        \sample_f2_wdata[66]\, sample_f2_wdata(65) => 
        \sample_f2_wdata[65]\, sample_f2_wdata(64) => 
        \sample_f2_wdata[64]\, sample_f2_wdata(63) => 
        \sample_f2_wdata[63]\, sample_f2_wdata(62) => 
        \sample_f2_wdata[62]\, sample_f2_wdata(61) => 
        \sample_f2_wdata[61]\, sample_f2_wdata(60) => 
        \sample_f2_wdata[60]\, sample_f2_wdata(59) => 
        \sample_f2_wdata[59]\, sample_f2_wdata(58) => 
        \sample_f2_wdata[58]\, sample_f2_wdata(57) => 
        \sample_f2_wdata[57]\, sample_f2_wdata(56) => 
        \sample_f2_wdata[56]\, sample_f2_wdata(55) => 
        \sample_f2_wdata[55]\, sample_f2_wdata(54) => 
        \sample_f2_wdata[54]\, sample_f2_wdata(53) => 
        \sample_f2_wdata[53]\, sample_f2_wdata(52) => 
        \sample_f2_wdata[52]\, sample_f2_wdata(51) => 
        \sample_f2_wdata[51]\, sample_f2_wdata(50) => 
        \sample_f2_wdata[50]\, sample_f2_wdata(49) => 
        \sample_f2_wdata[49]\, sample_f2_wdata(48) => 
        \sample_f2_wdata[48]\, sample_f2_wdata(47) => 
        \sample_f2_wdata[47]\, sample_f2_wdata(46) => 
        \sample_f2_wdata[46]\, sample_f2_wdata(45) => 
        \sample_f2_wdata[45]\, sample_f2_wdata(44) => 
        \sample_f2_wdata[44]\, sample_f2_wdata(43) => 
        \sample_f2_wdata[43]\, sample_f2_wdata(42) => 
        \sample_f2_wdata[42]\, sample_f2_wdata(41) => 
        \sample_f2_wdata[41]\, sample_f2_wdata(40) => 
        \sample_f2_wdata[40]\, sample_f2_wdata(39) => 
        \sample_f2_wdata[39]\, sample_f2_wdata(38) => 
        \sample_f2_wdata[38]\, sample_f2_wdata(37) => 
        \sample_f2_wdata[37]\, sample_f2_wdata(36) => 
        \sample_f2_wdata[36]\, sample_f2_wdata(35) => 
        \sample_f2_wdata[35]\, sample_f2_wdata(34) => 
        \sample_f2_wdata[34]\, sample_f2_wdata(33) => 
        \sample_f2_wdata[33]\, sample_f2_wdata(32) => 
        \sample_f2_wdata[32]\, sample_f2_wdata(31) => 
        \sample_f2_wdata[31]\, sample_f2_wdata(30) => 
        \sample_f2_wdata[30]\, sample_f2_wdata(29) => 
        \sample_f2_wdata[29]\, sample_f2_wdata(28) => 
        \sample_f2_wdata[28]\, sample_f2_wdata(27) => 
        \sample_f2_wdata[27]\, sample_f2_wdata(26) => 
        \sample_f2_wdata[26]\, sample_f2_wdata(25) => 
        \sample_f2_wdata[25]\, sample_f2_wdata(24) => 
        \sample_f2_wdata[24]\, sample_f2_wdata(23) => 
        \sample_f2_wdata[23]\, sample_f2_wdata(22) => 
        \sample_f2_wdata[22]\, sample_f2_wdata(21) => 
        \sample_f2_wdata[21]\, sample_f2_wdata(20) => 
        \sample_f2_wdata[20]\, sample_f2_wdata(19) => 
        \sample_f2_wdata[19]\, sample_f2_wdata(18) => 
        \sample_f2_wdata[18]\, sample_f2_wdata(17) => 
        \sample_f2_wdata[17]\, sample_f2_wdata(16) => 
        \sample_f2_wdata[16]\, sample_f2_wdata(15) => 
        \sample_f2_wdata[15]\, sample_f2_wdata(14) => 
        \sample_f2_wdata[14]\, sample_f2_wdata(13) => 
        \sample_f2_wdata[13]\, sample_f2_wdata(12) => 
        \sample_f2_wdata[12]\, sample_f2_wdata(11) => 
        \sample_f2_wdata[11]\, sample_f2_wdata(10) => 
        \sample_f2_wdata[10]\, sample_f2_wdata(9) => 
        \sample_f2_wdata[9]\, sample_f2_wdata(8) => 
        \sample_f2_wdata[8]\, sample_f2_wdata(7) => 
        \sample_f2_wdata[7]\, sample_f2_wdata(6) => 
        \sample_f2_wdata[6]\, sample_f2_wdata(5) => 
        \sample_f2_wdata[5]\, sample_f2_wdata(4) => 
        \sample_f2_wdata[4]\, sample_f2_wdata(3) => 
        \sample_f2_wdata[3]\, sample_f2_wdata(2) => 
        \sample_f2_wdata[2]\, sample_f2_wdata(1) => 
        \sample_f2_wdata[1]\, sample_f2_wdata(0) => 
        \sample_f2_wdata[0]\, sample_f0_val => sample_f0_val, 
        sample_f0_val_1 => sample_f0_val_1, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, sample_f2_val => 
        sample_f2_val, sample_f0_val_0 => sample_f0_val_0, 
        sample_out_0_sqmuxa_1 => sample_out_0_sqmuxa_1);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I38_Y : 
        AO13
      port map(A => N194_0, B => \sample_filter_v2_out[99]\, C
         => \sample_filter_v2_out[117]\, Y => N264_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I95_Y_0 : 
        XOR3
      port map(A => \sample_filter_v2_out[105]\, B => 
        \sample_filter_v2_out[123]\, C => N294_i, Y => 
        \sample_data_shaping_f2_f1_s[2]\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[33]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[33]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[33]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I53_Y : 
        OR2B
      port map(A => SUB_16x16_medium_area_I53_Y_0_0, B => 
        I53_un1_Y, Y => N278);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I56_Y : 
        AO1B
      port map(A => SUB_16x16_medium_area_I56_un1_Y_0, B => N278, 
        C => SUB_16x16_medium_area_I56_Y_1_0, Y => N268);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out_RNO[111]\ : 
        MX2B
      port map(A => \sample_filter_v2_out[111]\, B => 
        \sample_data_shaping_f1_f0_s_i[14]\, S => 
        data_shaping_SP0, Y => \sample_data_shaping_out_349[111]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I89_Y : 
        AO18
      port map(A => N268, B => \sample_filter_v2_out[136]\, C => 
        \sample_filter_v2_out[118]\, Y => N288_i);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[122]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_85[122]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[122]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[20]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[20]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[20]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I53_Y : 
        AO1B
      port map(A => SUB_16x16_medium_area_I53_un1_Y_0, B => 
        N181_0, C => SUB_16x16_medium_area_I53_Y_0, Y => N278_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I87_Y : 
        AO18
      port map(A => N258, B => \sample_filter_v2_out[132]\, C => 
        \sample_filter_v2_out[114]\, Y => N284_i);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out_RNO[96]\ : 
        MX2
      port map(A => \sample_filter_v2_out[96]\, B => 
        \sample_data_shaping_f2_f1_s[11]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_281[96]\);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[3]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[3]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[3]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I57_un1_Y_0 : 
        NOR2B
      port map(A => N229_0, B => N245_0, Y => 
        SUB_16x16_medium_area_I57_un1_Y_0_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I43_Y : 
        NOR2B
      port map(A => N187, B => N185, Y => N275);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[58]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[58]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[58]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I46_Y : 
        OR2A
      port map(A => \sample_filter_v2_out[143]\, B => 
        \sample_filter_v2_out[125]\, Y => N225_0);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[26]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[26]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[26]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[56]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[56]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[56]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I102_Y_0 : 
        AX1D
      port map(A => I78_un1_Y, B => N264_0, C => N197_0, Y => 
        \sample_data_shaping_f2_f1_s[9]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I21_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[138]\, B => 
        \sample_filter_v2_out[120]\, Y => N189);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[143]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[143]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[143]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I26_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[115]\, B => 
        \sample_filter_v2_out[97]\, Y => N199);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I88_un1_Y : 
        OA1
      port map(A => I78_un1_Y, B => N264_0, C => N197_0, Y => 
        I88_un1_Y);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out_RNO[107]\ : 
        AX1C
      port map(A => \sample_filter_v2_out[125]\, B => 
        data_shaping_SP1, C => \sample_filter_v2_out[107]\, Y => 
        \sample_data_shaping_out_17[107]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I85_Y : 
        AO1
      port map(A => N278_0, B => N275_0, C => N274, Y => N280);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[27]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[27]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[27]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I85_un1_Y : 
        NOR2B
      port map(A => N278, B => N275, Y => I85_un1_Y);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[136]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[136]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[136]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I39_Y : 
        XA1A
      port map(A => \sample_filter_v2_out[118]\, B => 
        \sample_filter_v2_out[136]\, C => N195, Y => N265);
    
    lpp_waveform_1 : lpp_waveform
      port map(status_full_ack(3) => status_full_ack(3), 
        status_full_ack(2) => status_full_ack(2), 
        status_full_ack(1) => status_full_ack(1), 
        status_full_ack(0) => status_full_ack(0), hburst_c(2) => 
        hburst_c(2), hburst_c(1) => hburst_c(1), hburst_c(0) => 
        hburst_c(0), htrans_c(1) => htrans_c(1), htrans_c(0) => 
        htrans_c(0), hsize_c(1) => hsize_c(1), hsize_c(0) => 
        hsize_c(0), AHB_Master_In_c_5 => AHB_Master_In_c_5, 
        AHB_Master_In_c_4 => AHB_Master_In_c_4, AHB_Master_In_c_0
         => AHB_Master_In_c_0, AHB_Master_In_c_3 => 
        AHB_Master_In_c_3, haddr_c(31) => haddr_c(31), 
        haddr_c(30) => haddr_c(30), haddr_c(29) => haddr_c(29), 
        haddr_c(28) => haddr_c(28), haddr_c(27) => haddr_c(27), 
        haddr_c(26) => haddr_c(26), haddr_c(25) => haddr_c(25), 
        haddr_c(24) => haddr_c(24), haddr_c(23) => haddr_c(23), 
        haddr_c(22) => haddr_c(22), haddr_c(21) => haddr_c(21), 
        haddr_c(20) => haddr_c(20), haddr_c(19) => haddr_c(19), 
        haddr_c(18) => haddr_c(18), haddr_c(17) => haddr_c(17), 
        haddr_c(16) => haddr_c(16), haddr_c(15) => haddr_c(15), 
        haddr_c(14) => haddr_c(14), haddr_c(13) => haddr_c(13), 
        haddr_c(12) => haddr_c(12), haddr_c(11) => haddr_c(11), 
        haddr_c(10) => haddr_c(10), haddr_c(9) => haddr_c(9), 
        haddr_c(8) => haddr_c(8), haddr_c(7) => haddr_c(7), 
        haddr_c(6) => haddr_c(6), haddr_c(5) => haddr_c(5), 
        haddr_c(4) => haddr_c(4), haddr_c(3) => haddr_c(3), 
        haddr_c(2) => haddr_c(2), haddr_c(1) => haddr_c(1), 
        haddr_c(0) => haddr_c(0), nb_burst_available(10) => 
        nb_burst_available(10), nb_burst_available(9) => 
        nb_burst_available(9), nb_burst_available(8) => 
        nb_burst_available(8), nb_burst_available(7) => 
        nb_burst_available(7), nb_burst_available(6) => 
        nb_burst_available(6), nb_burst_available(5) => 
        nb_burst_available(5), nb_burst_available(4) => 
        nb_burst_available(4), nb_burst_available(3) => 
        nb_burst_available(3), nb_burst_available(2) => 
        nb_burst_available(2), nb_burst_available(1) => 
        nb_burst_available(1), nb_burst_available(0) => 
        nb_burst_available(0), status_full_err(3) => 
        status_full_err(3), status_full_err(2) => 
        status_full_err(2), status_full_err(1) => 
        status_full_err(1), status_full_err(0) => 
        status_full_err(0), status_full(3) => status_full(3), 
        status_full(2) => status_full(2), status_full(1) => 
        status_full(1), status_full(0) => status_full(0), 
        addr_data_f3(31) => addr_data_f3(31), addr_data_f3(30)
         => addr_data_f3(30), addr_data_f3(29) => 
        addr_data_f3(29), addr_data_f3(28) => addr_data_f3(28), 
        addr_data_f3(27) => addr_data_f3(27), addr_data_f3(26)
         => addr_data_f3(26), addr_data_f3(25) => 
        addr_data_f3(25), addr_data_f3(24) => addr_data_f3(24), 
        addr_data_f3(23) => addr_data_f3(23), addr_data_f3(22)
         => addr_data_f3(22), addr_data_f3(21) => 
        addr_data_f3(21), addr_data_f3(20) => addr_data_f3(20), 
        addr_data_f3(19) => addr_data_f3(19), addr_data_f3(18)
         => addr_data_f3(18), addr_data_f3(17) => 
        addr_data_f3(17), addr_data_f3(16) => addr_data_f3(16), 
        addr_data_f3(15) => addr_data_f3(15), addr_data_f3(14)
         => addr_data_f3(14), addr_data_f3(13) => 
        addr_data_f3(13), addr_data_f3(12) => addr_data_f3(12), 
        addr_data_f3(11) => addr_data_f3(11), addr_data_f3(10)
         => addr_data_f3(10), addr_data_f3(9) => addr_data_f3(9), 
        addr_data_f3(8) => addr_data_f3(8), addr_data_f3(7) => 
        addr_data_f3(7), addr_data_f3(6) => addr_data_f3(6), 
        addr_data_f3(5) => addr_data_f3(5), addr_data_f3(4) => 
        addr_data_f3(4), addr_data_f3(3) => addr_data_f3(3), 
        addr_data_f3(2) => addr_data_f3(2), addr_data_f3(1) => 
        addr_data_f3(1), addr_data_f3(0) => addr_data_f3(0), 
        addr_data_f2(31) => addr_data_f2(31), addr_data_f2(30)
         => addr_data_f2(30), addr_data_f2(29) => 
        addr_data_f2(29), addr_data_f2(28) => addr_data_f2(28), 
        addr_data_f2(27) => addr_data_f2(27), addr_data_f2(26)
         => addr_data_f2(26), addr_data_f2(25) => 
        addr_data_f2(25), addr_data_f2(24) => addr_data_f2(24), 
        addr_data_f2(23) => addr_data_f2(23), addr_data_f2(22)
         => addr_data_f2(22), addr_data_f2(21) => 
        addr_data_f2(21), addr_data_f2(20) => addr_data_f2(20), 
        addr_data_f2(19) => addr_data_f2(19), addr_data_f2(18)
         => addr_data_f2(18), addr_data_f2(17) => 
        addr_data_f2(17), addr_data_f2(16) => addr_data_f2(16), 
        addr_data_f2(15) => addr_data_f2(15), addr_data_f2(14)
         => addr_data_f2(14), addr_data_f2(13) => 
        addr_data_f2(13), addr_data_f2(12) => addr_data_f2(12), 
        addr_data_f2(11) => addr_data_f2(11), addr_data_f2(10)
         => addr_data_f2(10), addr_data_f2(9) => addr_data_f2(9), 
        addr_data_f2(8) => addr_data_f2(8), addr_data_f2(7) => 
        addr_data_f2(7), addr_data_f2(6) => addr_data_f2(6), 
        addr_data_f2(5) => addr_data_f2(5), addr_data_f2(4) => 
        addr_data_f2(4), addr_data_f2(3) => addr_data_f2(3), 
        addr_data_f2(2) => addr_data_f2(2), addr_data_f2(1) => 
        addr_data_f2(1), addr_data_f2(0) => addr_data_f2(0), 
        addr_data_f1(31) => addr_data_f1(31), addr_data_f1(30)
         => addr_data_f1(30), addr_data_f1(29) => 
        addr_data_f1(29), addr_data_f1(28) => addr_data_f1(28), 
        addr_data_f1(27) => addr_data_f1(27), addr_data_f1(26)
         => addr_data_f1(26), addr_data_f1(25) => 
        addr_data_f1(25), addr_data_f1(24) => addr_data_f1(24), 
        addr_data_f1(23) => addr_data_f1(23), addr_data_f1(22)
         => addr_data_f1(22), addr_data_f1(21) => 
        addr_data_f1(21), addr_data_f1(20) => addr_data_f1(20), 
        addr_data_f1(19) => addr_data_f1(19), addr_data_f1(18)
         => addr_data_f1(18), addr_data_f1(17) => 
        addr_data_f1(17), addr_data_f1(16) => addr_data_f1(16), 
        addr_data_f1(15) => addr_data_f1(15), addr_data_f1(14)
         => addr_data_f1(14), addr_data_f1(13) => 
        addr_data_f1(13), addr_data_f1(12) => addr_data_f1(12), 
        addr_data_f1(11) => addr_data_f1(11), addr_data_f1(10)
         => addr_data_f1(10), addr_data_f1(9) => addr_data_f1(9), 
        addr_data_f1(8) => addr_data_f1(8), addr_data_f1(7) => 
        addr_data_f1(7), addr_data_f1(6) => addr_data_f1(6), 
        addr_data_f1(5) => addr_data_f1(5), addr_data_f1(4) => 
        addr_data_f1(4), addr_data_f1(3) => addr_data_f1(3), 
        addr_data_f1(2) => addr_data_f1(2), addr_data_f1(1) => 
        addr_data_f1(1), addr_data_f1(0) => addr_data_f1(0), 
        addr_data_f0(31) => addr_data_f0(31), addr_data_f0(30)
         => addr_data_f0(30), addr_data_f0(29) => 
        addr_data_f0(29), addr_data_f0(28) => addr_data_f0(28), 
        addr_data_f0(27) => addr_data_f0(27), addr_data_f0(26)
         => addr_data_f0(26), addr_data_f0(25) => 
        addr_data_f0(25), addr_data_f0(24) => addr_data_f0(24), 
        addr_data_f0(23) => addr_data_f0(23), addr_data_f0(22)
         => addr_data_f0(22), addr_data_f0(21) => 
        addr_data_f0(21), addr_data_f0(20) => addr_data_f0(20), 
        addr_data_f0(19) => addr_data_f0(19), addr_data_f0(18)
         => addr_data_f0(18), addr_data_f0(17) => 
        addr_data_f0(17), addr_data_f0(16) => addr_data_f0(16), 
        addr_data_f0(15) => addr_data_f0(15), addr_data_f0(14)
         => addr_data_f0(14), addr_data_f0(13) => 
        addr_data_f0(13), addr_data_f0(12) => addr_data_f0(12), 
        addr_data_f0(11) => addr_data_f0(11), addr_data_f0(10)
         => addr_data_f0(10), addr_data_f0(9) => addr_data_f0(9), 
        addr_data_f0(8) => addr_data_f0(8), addr_data_f0(7) => 
        addr_data_f0(7), addr_data_f0(6) => addr_data_f0(6), 
        addr_data_f0(5) => addr_data_f0(5), addr_data_f0(4) => 
        addr_data_f0(4), addr_data_f0(3) => addr_data_f0(3), 
        addr_data_f0(2) => addr_data_f0(2), addr_data_f0(1) => 
        addr_data_f0(1), addr_data_f0(0) => addr_data_f0(0), 
        hwdata_c(31) => hwdata_c(31), hwdata_c(30) => 
        hwdata_c(30), hwdata_c(29) => hwdata_c(29), hwdata_c(28)
         => hwdata_c(28), hwdata_c(27) => hwdata_c(27), 
        hwdata_c(26) => hwdata_c(26), hwdata_c(25) => 
        hwdata_c(25), hwdata_c(24) => hwdata_c(24), hwdata_c(23)
         => hwdata_c(23), hwdata_c(22) => hwdata_c(22), 
        hwdata_c(21) => hwdata_c(21), hwdata_c(20) => 
        hwdata_c(20), hwdata_c(19) => hwdata_c(19), hwdata_c(18)
         => hwdata_c(18), hwdata_c(17) => hwdata_c(17), 
        hwdata_c(16) => hwdata_c(16), hwdata_c(15) => 
        hwdata_c(15), hwdata_c(14) => hwdata_c(14), hwdata_c(13)
         => hwdata_c(13), hwdata_c(12) => hwdata_c(12), 
        hwdata_c(11) => hwdata_c(11), hwdata_c(10) => 
        hwdata_c(10), hwdata_c(9) => hwdata_c(9), hwdata_c(8) => 
        hwdata_c(8), hwdata_c(7) => hwdata_c(7), hwdata_c(6) => 
        hwdata_c(6), hwdata_c(5) => hwdata_c(5), hwdata_c(4) => 
        hwdata_c(4), hwdata_c(3) => hwdata_c(3), hwdata_c(2) => 
        hwdata_c(2), hwdata_c(1) => hwdata_c(1), hwdata_c(0) => 
        hwdata_c(0), status_new_err(3) => status_new_err(3), 
        status_new_err(2) => status_new_err(2), status_new_err(1)
         => status_new_err(1), status_new_err(0) => 
        status_new_err(0), sample_f3_wdata(95) => 
        \sample_f3_wdata[95]\, sample_f3_wdata(94) => 
        \sample_f3_wdata[94]\, sample_f3_wdata(93) => 
        \sample_f3_wdata[93]\, sample_f3_wdata(92) => 
        \sample_f3_wdata[92]\, sample_f3_wdata(91) => 
        \sample_f3_wdata[91]\, sample_f3_wdata(90) => 
        \sample_f3_wdata[90]\, sample_f3_wdata(89) => 
        \sample_f3_wdata[89]\, sample_f3_wdata(88) => 
        \sample_f3_wdata[88]\, sample_f3_wdata(87) => 
        \sample_f3_wdata[87]\, sample_f3_wdata(86) => 
        \sample_f3_wdata[86]\, sample_f3_wdata(85) => 
        \sample_f3_wdata[85]\, sample_f3_wdata(84) => 
        \sample_f3_wdata[84]\, sample_f3_wdata(83) => 
        \sample_f3_wdata[83]\, sample_f3_wdata(82) => 
        \sample_f3_wdata[82]\, sample_f3_wdata(81) => 
        \sample_f3_wdata[81]\, sample_f3_wdata(80) => 
        \sample_f3_wdata[80]\, sample_f3_wdata(79) => 
        \sample_f3_wdata[79]\, sample_f3_wdata(78) => 
        \sample_f3_wdata[78]\, sample_f3_wdata(77) => 
        \sample_f3_wdata[77]\, sample_f3_wdata(76) => 
        \sample_f3_wdata[76]\, sample_f3_wdata(75) => 
        \sample_f3_wdata[75]\, sample_f3_wdata(74) => 
        \sample_f3_wdata[74]\, sample_f3_wdata(73) => 
        \sample_f3_wdata[73]\, sample_f3_wdata(72) => 
        \sample_f3_wdata[72]\, sample_f3_wdata(71) => 
        \sample_f3_wdata[71]\, sample_f3_wdata(70) => 
        \sample_f3_wdata[70]\, sample_f3_wdata(69) => 
        \sample_f3_wdata[69]\, sample_f3_wdata(68) => 
        \sample_f3_wdata[68]\, sample_f3_wdata(67) => 
        \sample_f3_wdata[67]\, sample_f3_wdata(66) => 
        \sample_f3_wdata[66]\, sample_f3_wdata(65) => 
        \sample_f3_wdata[65]\, sample_f3_wdata(64) => 
        \sample_f3_wdata[64]\, sample_f3_wdata(63) => 
        \sample_f3_wdata[63]\, sample_f3_wdata(62) => 
        \sample_f3_wdata[62]\, sample_f3_wdata(61) => 
        \sample_f3_wdata[61]\, sample_f3_wdata(60) => 
        \sample_f3_wdata[60]\, sample_f3_wdata(59) => 
        \sample_f3_wdata[59]\, sample_f3_wdata(58) => 
        \sample_f3_wdata[58]\, sample_f3_wdata(57) => 
        \sample_f3_wdata[57]\, sample_f3_wdata(56) => 
        \sample_f3_wdata[56]\, sample_f3_wdata(55) => 
        \sample_f3_wdata[55]\, sample_f3_wdata(54) => 
        \sample_f3_wdata[54]\, sample_f3_wdata(53) => 
        \sample_f3_wdata[53]\, sample_f3_wdata(52) => 
        \sample_f3_wdata[52]\, sample_f3_wdata(51) => 
        \sample_f3_wdata[51]\, sample_f3_wdata(50) => 
        \sample_f3_wdata[50]\, sample_f3_wdata(49) => 
        \sample_f3_wdata[49]\, sample_f3_wdata(48) => 
        \sample_f3_wdata[48]\, sample_f3_wdata(47) => 
        \sample_f3_wdata[47]\, sample_f3_wdata(46) => 
        \sample_f3_wdata[46]\, sample_f3_wdata(45) => 
        \sample_f3_wdata[45]\, sample_f3_wdata(44) => 
        \sample_f3_wdata[44]\, sample_f3_wdata(43) => 
        \sample_f3_wdata[43]\, sample_f3_wdata(42) => 
        \sample_f3_wdata[42]\, sample_f3_wdata(41) => 
        \sample_f3_wdata[41]\, sample_f3_wdata(40) => 
        \sample_f3_wdata[40]\, sample_f3_wdata(39) => 
        \sample_f3_wdata[39]\, sample_f3_wdata(38) => 
        \sample_f3_wdata[38]\, sample_f3_wdata(37) => 
        \sample_f3_wdata[37]\, sample_f3_wdata(36) => 
        \sample_f3_wdata[36]\, sample_f3_wdata(35) => 
        \sample_f3_wdata[35]\, sample_f3_wdata(34) => 
        \sample_f3_wdata[34]\, sample_f3_wdata(33) => 
        \sample_f3_wdata[33]\, sample_f3_wdata(32) => 
        \sample_f3_wdata[32]\, sample_f3_wdata(31) => 
        \sample_f3_wdata[31]\, sample_f3_wdata(30) => 
        \sample_f3_wdata[30]\, sample_f3_wdata(29) => 
        \sample_f3_wdata[29]\, sample_f3_wdata(28) => 
        \sample_f3_wdata[28]\, sample_f3_wdata(27) => 
        \sample_f3_wdata[27]\, sample_f3_wdata(26) => 
        \sample_f3_wdata[26]\, sample_f3_wdata(25) => 
        \sample_f3_wdata[25]\, sample_f3_wdata(24) => 
        \sample_f3_wdata[24]\, sample_f3_wdata(23) => 
        \sample_f3_wdata[23]\, sample_f3_wdata(22) => 
        \sample_f3_wdata[22]\, sample_f3_wdata(21) => 
        \sample_f3_wdata[21]\, sample_f3_wdata(20) => 
        \sample_f3_wdata[20]\, sample_f3_wdata(19) => 
        \sample_f3_wdata[19]\, sample_f3_wdata(18) => 
        \sample_f3_wdata[18]\, sample_f3_wdata(17) => 
        \sample_f3_wdata[17]\, sample_f3_wdata(16) => 
        \sample_f3_wdata[16]\, sample_f3_wdata(15) => 
        \sample_f3_wdata[15]\, sample_f3_wdata(14) => 
        \sample_f3_wdata[14]\, sample_f3_wdata(13) => 
        \sample_f3_wdata[13]\, sample_f3_wdata(12) => 
        \sample_f3_wdata[12]\, sample_f3_wdata(11) => 
        \sample_f3_wdata[11]\, sample_f3_wdata(10) => 
        \sample_f3_wdata[10]\, sample_f3_wdata(9) => 
        \sample_f3_wdata[9]\, sample_f3_wdata(8) => 
        \sample_f3_wdata[8]\, sample_f3_wdata(7) => 
        \sample_f3_wdata[7]\, sample_f3_wdata(6) => 
        \sample_f3_wdata[6]\, sample_f3_wdata(5) => 
        \sample_f3_wdata[5]\, sample_f3_wdata(4) => 
        \sample_f3_wdata[4]\, sample_f3_wdata(3) => 
        \sample_f3_wdata[3]\, sample_f3_wdata(2) => 
        \sample_f3_wdata[2]\, sample_f3_wdata(1) => 
        \sample_f3_wdata[1]\, sample_f3_wdata(0) => 
        \sample_f3_wdata[0]\, sample_f2_wdata(95) => 
        \sample_f2_wdata[95]\, sample_f2_wdata(94) => 
        \sample_f2_wdata[94]\, sample_f2_wdata(93) => 
        \sample_f2_wdata[93]\, sample_f2_wdata(92) => 
        \sample_f2_wdata[92]\, sample_f2_wdata(91) => 
        \sample_f2_wdata[91]\, sample_f2_wdata(90) => 
        \sample_f2_wdata[90]\, sample_f2_wdata(89) => 
        \sample_f2_wdata[89]\, sample_f2_wdata(88) => 
        \sample_f2_wdata[88]\, sample_f2_wdata(87) => 
        \sample_f2_wdata[87]\, sample_f2_wdata(86) => 
        \sample_f2_wdata[86]\, sample_f2_wdata(85) => 
        \sample_f2_wdata[85]\, sample_f2_wdata(84) => 
        \sample_f2_wdata[84]\, sample_f2_wdata(83) => 
        \sample_f2_wdata[83]\, sample_f2_wdata(82) => 
        \sample_f2_wdata[82]\, sample_f2_wdata(81) => 
        \sample_f2_wdata[81]\, sample_f2_wdata(80) => 
        \sample_f2_wdata[80]\, sample_f2_wdata(79) => 
        \sample_f2_wdata[79]\, sample_f2_wdata(78) => 
        \sample_f2_wdata[78]\, sample_f2_wdata(77) => 
        \sample_f2_wdata[77]\, sample_f2_wdata(76) => 
        \sample_f2_wdata[76]\, sample_f2_wdata(75) => 
        \sample_f2_wdata[75]\, sample_f2_wdata(74) => 
        \sample_f2_wdata[74]\, sample_f2_wdata(73) => 
        \sample_f2_wdata[73]\, sample_f2_wdata(72) => 
        \sample_f2_wdata[72]\, sample_f2_wdata(71) => 
        \sample_f2_wdata[71]\, sample_f2_wdata(70) => 
        \sample_f2_wdata[70]\, sample_f2_wdata(69) => 
        \sample_f2_wdata[69]\, sample_f2_wdata(68) => 
        \sample_f2_wdata[68]\, sample_f2_wdata(67) => 
        \sample_f2_wdata[67]\, sample_f2_wdata(66) => 
        \sample_f2_wdata[66]\, sample_f2_wdata(65) => 
        \sample_f2_wdata[65]\, sample_f2_wdata(64) => 
        \sample_f2_wdata[64]\, sample_f2_wdata(63) => 
        \sample_f2_wdata[63]\, sample_f2_wdata(62) => 
        \sample_f2_wdata[62]\, sample_f2_wdata(61) => 
        \sample_f2_wdata[61]\, sample_f2_wdata(60) => 
        \sample_f2_wdata[60]\, sample_f2_wdata(59) => 
        \sample_f2_wdata[59]\, sample_f2_wdata(58) => 
        \sample_f2_wdata[58]\, sample_f2_wdata(57) => 
        \sample_f2_wdata[57]\, sample_f2_wdata(56) => 
        \sample_f2_wdata[56]\, sample_f2_wdata(55) => 
        \sample_f2_wdata[55]\, sample_f2_wdata(54) => 
        \sample_f2_wdata[54]\, sample_f2_wdata(53) => 
        \sample_f2_wdata[53]\, sample_f2_wdata(52) => 
        \sample_f2_wdata[52]\, sample_f2_wdata(51) => 
        \sample_f2_wdata[51]\, sample_f2_wdata(50) => 
        \sample_f2_wdata[50]\, sample_f2_wdata(49) => 
        \sample_f2_wdata[49]\, sample_f2_wdata(48) => 
        \sample_f2_wdata[48]\, sample_f2_wdata(47) => 
        \sample_f2_wdata[47]\, sample_f2_wdata(46) => 
        \sample_f2_wdata[46]\, sample_f2_wdata(45) => 
        \sample_f2_wdata[45]\, sample_f2_wdata(44) => 
        \sample_f2_wdata[44]\, sample_f2_wdata(43) => 
        \sample_f2_wdata[43]\, sample_f2_wdata(42) => 
        \sample_f2_wdata[42]\, sample_f2_wdata(41) => 
        \sample_f2_wdata[41]\, sample_f2_wdata(40) => 
        \sample_f2_wdata[40]\, sample_f2_wdata(39) => 
        \sample_f2_wdata[39]\, sample_f2_wdata(38) => 
        \sample_f2_wdata[38]\, sample_f2_wdata(37) => 
        \sample_f2_wdata[37]\, sample_f2_wdata(36) => 
        \sample_f2_wdata[36]\, sample_f2_wdata(35) => 
        \sample_f2_wdata[35]\, sample_f2_wdata(34) => 
        \sample_f2_wdata[34]\, sample_f2_wdata(33) => 
        \sample_f2_wdata[33]\, sample_f2_wdata(32) => 
        \sample_f2_wdata[32]\, sample_f2_wdata(31) => 
        \sample_f2_wdata[31]\, sample_f2_wdata(30) => 
        \sample_f2_wdata[30]\, sample_f2_wdata(29) => 
        \sample_f2_wdata[29]\, sample_f2_wdata(28) => 
        \sample_f2_wdata[28]\, sample_f2_wdata(27) => 
        \sample_f2_wdata[27]\, sample_f2_wdata(26) => 
        \sample_f2_wdata[26]\, sample_f2_wdata(25) => 
        \sample_f2_wdata[25]\, sample_f2_wdata(24) => 
        \sample_f2_wdata[24]\, sample_f2_wdata(23) => 
        \sample_f2_wdata[23]\, sample_f2_wdata(22) => 
        \sample_f2_wdata[22]\, sample_f2_wdata(21) => 
        \sample_f2_wdata[21]\, sample_f2_wdata(20) => 
        \sample_f2_wdata[20]\, sample_f2_wdata(19) => 
        \sample_f2_wdata[19]\, sample_f2_wdata(18) => 
        \sample_f2_wdata[18]\, sample_f2_wdata(17) => 
        \sample_f2_wdata[17]\, sample_f2_wdata(16) => 
        \sample_f2_wdata[16]\, sample_f2_wdata(15) => 
        \sample_f2_wdata[15]\, sample_f2_wdata(14) => 
        \sample_f2_wdata[14]\, sample_f2_wdata(13) => 
        \sample_f2_wdata[13]\, sample_f2_wdata(12) => 
        \sample_f2_wdata[12]\, sample_f2_wdata(11) => 
        \sample_f2_wdata[11]\, sample_f2_wdata(10) => 
        \sample_f2_wdata[10]\, sample_f2_wdata(9) => 
        \sample_f2_wdata[9]\, sample_f2_wdata(8) => 
        \sample_f2_wdata[8]\, sample_f2_wdata(7) => 
        \sample_f2_wdata[7]\, sample_f2_wdata(6) => 
        \sample_f2_wdata[6]\, sample_f2_wdata(5) => 
        \sample_f2_wdata[5]\, sample_f2_wdata(4) => 
        \sample_f2_wdata[4]\, sample_f2_wdata(3) => 
        \sample_f2_wdata[3]\, sample_f2_wdata(2) => 
        \sample_f2_wdata[2]\, sample_f2_wdata(1) => 
        \sample_f2_wdata[1]\, sample_f2_wdata(0) => 
        \sample_f2_wdata[0]\, sample_f1_15 => \sample_f1[63]\, 
        sample_f1_47 => \sample_f1[95]\, sample_f1_14 => 
        \sample_f1[62]\, sample_f1_46 => \sample_f1[94]\, 
        sample_f1_13 => \sample_f1[61]\, sample_f1_45 => 
        \sample_f1[93]\, sample_f1_12 => \sample_f1[60]\, 
        sample_f1_44 => \sample_f1[92]\, sample_f1_60 => 
        \sample_f1[108]\, sample_f1_59 => \sample_f1[107]\, 
        sample_f1_58 => \sample_f1[106]\, sample_f1_57 => 
        \sample_f1[105]\, sample_f1_56 => \sample_f1[104]\, 
        sample_f1_55 => \sample_f1[103]\, sample_f1_54 => 
        \sample_f1[102]\, sample_f1_53 => \sample_f1[101]\, 
        sample_f1_52 => \sample_f1[100]\, sample_f1_51 => 
        \sample_f1[99]\, sample_f1_50 => \sample_f1[98]\, 
        sample_f1_49 => \sample_f1[97]\, sample_f1_48 => 
        \sample_f1[96]\, sample_f1_4 => \sample_f1[52]\, 
        sample_f1_36 => \sample_f1[84]\, sample_f1_3 => 
        \sample_f1[51]\, sample_f1_35 => \sample_f1[83]\, 
        sample_f1_2 => \sample_f1[50]\, sample_f1_34 => 
        \sample_f1[82]\, sample_f1_1 => \sample_f1[49]\, 
        sample_f1_33 => \sample_f1[81]\, sample_f1_0 => 
        \sample_f1[48]\, sample_f1_32 => \sample_f1[80]\, 
        sample_f1_63 => \sample_f1[111]\, sample_f1_62 => 
        \sample_f1[110]\, sample_f1_61 => \sample_f1[109]\, 
        sample_f1_11 => \sample_f1[59]\, sample_f1_43 => 
        \sample_f1[91]\, sample_f1_10 => \sample_f1[58]\, 
        sample_f1_42 => \sample_f1[90]\, sample_f1_9 => 
        \sample_f1[57]\, sample_f1_41 => \sample_f1[89]\, 
        sample_f1_8 => \sample_f1[56]\, sample_f1_40 => 
        \sample_f1[88]\, sample_f1_7 => \sample_f1[55]\, 
        sample_f1_39 => \sample_f1[87]\, sample_f1_6 => 
        \sample_f1[54]\, sample_f1_38 => \sample_f1[86]\, 
        sample_f1_5 => \sample_f1[53]\, sample_f1_37 => 
        \sample_f1[85]\, sample_f1_wdata_0 => 
        \sample_f1_wdata[0]\, sample_f1_wdata_1 => 
        \sample_f1_wdata[1]\, sample_f1_wdata_2 => 
        \sample_f1_wdata[2]\, sample_f1_wdata_3 => 
        \sample_f1_wdata[3]\, sample_f1_wdata_4 => 
        \sample_f1_wdata[4]\, sample_f1_wdata_5 => 
        \sample_f1_wdata[5]\, sample_f1_wdata_6 => 
        \sample_f1_wdata[6]\, sample_f1_wdata_7 => 
        \sample_f1_wdata[7]\, sample_f1_wdata_8 => 
        \sample_f1_wdata[8]\, sample_f1_wdata_9 => 
        \sample_f1_wdata[9]\, sample_f1_wdata_10 => 
        \sample_f1_wdata[10]\, sample_f1_wdata_11 => 
        \sample_f1_wdata[11]\, sample_f1_wdata_12 => 
        \sample_f1_wdata[12]\, sample_f1_wdata_13 => 
        \sample_f1_wdata[13]\, sample_f1_wdata_14 => 
        \sample_f1_wdata[14]\, sample_f1_wdata_15 => 
        \sample_f1_wdata[15]\, sample_f1_wdata_48 => 
        \sample_f1_wdata[48]\, sample_f1_wdata_49 => 
        \sample_f1_wdata[49]\, sample_f1_wdata_50 => 
        \sample_f1_wdata[50]\, sample_f1_wdata_51 => 
        \sample_f1_wdata[51]\, sample_f1_wdata_52 => 
        \sample_f1_wdata[52]\, sample_f1_wdata_53 => 
        \sample_f1_wdata[53]\, sample_f1_wdata_54 => 
        \sample_f1_wdata[54]\, sample_f1_wdata_55 => 
        \sample_f1_wdata[55]\, sample_f1_wdata_56 => 
        \sample_f1_wdata[56]\, sample_f1_wdata_57 => 
        \sample_f1_wdata[57]\, sample_f1_wdata_58 => 
        \sample_f1_wdata[58]\, sample_f1_wdata_59 => 
        \sample_f1_wdata[59]\, sample_f1_wdata_60 => 
        \sample_f1_wdata[60]\, sample_f1_wdata_61 => 
        \sample_f1_wdata[61]\, sample_f1_wdata_62 => 
        \sample_f1_wdata[62]\, sample_f1_wdata_63 => 
        \sample_f1_wdata[63]\, sample_f1_wdata_64 => 
        \sample_f1_wdata[64]\, sample_f1_wdata_65 => 
        \sample_f1_wdata[65]\, sample_f1_wdata_66 => 
        \sample_f1_wdata[66]\, sample_f1_wdata_67 => 
        \sample_f1_wdata[67]\, sample_f1_wdata_68 => 
        \sample_f1_wdata[68]\, sample_f1_wdata_69 => 
        \sample_f1_wdata[69]\, sample_f1_wdata_70 => 
        \sample_f1_wdata[70]\, sample_f1_wdata_71 => 
        \sample_f1_wdata[71]\, sample_f1_wdata_72 => 
        \sample_f1_wdata[72]\, sample_f1_wdata_73 => 
        \sample_f1_wdata[73]\, sample_f1_wdata_74 => 
        \sample_f1_wdata[74]\, sample_f1_wdata_75 => 
        \sample_f1_wdata[75]\, sample_f1_wdata_76 => 
        \sample_f1_wdata[76]\, sample_f1_wdata_77 => 
        \sample_f1_wdata[77]\, sample_f1_wdata_78 => 
        \sample_f1_wdata[78]\, sample_f1_wdata_79 => 
        \sample_f1_wdata[79]\, sample_f1_wdata_80 => 
        \sample_f1_wdata[80]\, sample_f1_wdata_81 => 
        \sample_f1_wdata[81]\, sample_f1_wdata_82 => 
        \sample_f1_wdata[82]\, sample_f1_wdata_83 => 
        \sample_f1_wdata[83]\, sample_f1_wdata_84 => 
        \sample_f1_wdata[84]\, sample_f1_wdata_85 => 
        \sample_f1_wdata[85]\, sample_f1_wdata_86 => 
        \sample_f1_wdata[86]\, sample_f1_wdata_87 => 
        \sample_f1_wdata[87]\, sample_f1_wdata_88 => 
        \sample_f1_wdata[88]\, sample_f1_wdata_89 => 
        \sample_f1_wdata[89]\, sample_f1_wdata_90 => 
        \sample_f1_wdata[90]\, sample_f1_wdata_91 => 
        \sample_f1_wdata[91]\, sample_f1_wdata_92 => 
        \sample_f1_wdata[92]\, sample_f1_wdata_93 => 
        \sample_f1_wdata[93]\, sample_f1_wdata_94 => 
        \sample_f1_wdata[94]\, sample_f1_wdata_95 => 
        \sample_f1_wdata[95]\, sample_f0_15 => \sample_f0[63]\, 
        sample_f0_47 => \sample_f0[95]\, sample_f0_14 => 
        \sample_f0[62]\, sample_f0_46 => \sample_f0[94]\, 
        sample_f0_13 => \sample_f0[61]\, sample_f0_45 => 
        \sample_f0[93]\, sample_f0_12 => \sample_f0[60]\, 
        sample_f0_44 => \sample_f0[92]\, sample_f0_60 => 
        \sample_f0[108]\, sample_f0_59 => \sample_f0[107]\, 
        sample_f0_58 => \sample_f0[106]\, sample_f0_57 => 
        \sample_f0[105]\, sample_f0_56 => \sample_f0[104]\, 
        sample_f0_55 => \sample_f0[103]\, sample_f0_54 => 
        \sample_f0[102]\, sample_f0_53 => \sample_f0[101]\, 
        sample_f0_52 => \sample_f0[100]\, sample_f0_51 => 
        \sample_f0[99]\, sample_f0_50 => \sample_f0[98]\, 
        sample_f0_49 => \sample_f0[97]\, sample_f0_48 => 
        \sample_f0[96]\, sample_f0_4 => \sample_f0[52]\, 
        sample_f0_36 => \sample_f0[84]\, sample_f0_3 => 
        \sample_f0[51]\, sample_f0_35 => \sample_f0[83]\, 
        sample_f0_2 => \sample_f0[50]\, sample_f0_34 => 
        \sample_f0[82]\, sample_f0_1 => \sample_f0[49]\, 
        sample_f0_33 => \sample_f0[81]\, sample_f0_0 => 
        \sample_f0[48]\, sample_f0_32 => \sample_f0[80]\, 
        sample_f0_63 => \sample_f0[111]\, sample_f0_62 => 
        \sample_f0[110]\, sample_f0_61 => \sample_f0[109]\, 
        sample_f0_11 => \sample_f0[59]\, sample_f0_43 => 
        \sample_f0[91]\, sample_f0_10 => \sample_f0[58]\, 
        sample_f0_42 => \sample_f0[90]\, sample_f0_9 => 
        \sample_f0[57]\, sample_f0_41 => \sample_f0[89]\, 
        sample_f0_8 => \sample_f0[56]\, sample_f0_40 => 
        \sample_f0[88]\, sample_f0_7 => \sample_f0[55]\, 
        sample_f0_39 => \sample_f0[87]\, sample_f0_6 => 
        \sample_f0[54]\, sample_f0_38 => \sample_f0[86]\, 
        sample_f0_5 => \sample_f0[53]\, sample_f0_37 => 
        \sample_f0[85]\, sample_f0_wdata_0 => 
        \sample_f0_wdata[0]\, sample_f0_wdata_1 => 
        \sample_f0_wdata[1]\, sample_f0_wdata_2 => 
        \sample_f0_wdata[2]\, sample_f0_wdata_3 => 
        \sample_f0_wdata[3]\, sample_f0_wdata_4 => 
        \sample_f0_wdata[4]\, sample_f0_wdata_5 => 
        \sample_f0_wdata[5]\, sample_f0_wdata_6 => 
        \sample_f0_wdata[6]\, sample_f0_wdata_7 => 
        \sample_f0_wdata[7]\, sample_f0_wdata_8 => 
        \sample_f0_wdata[8]\, sample_f0_wdata_9 => 
        \sample_f0_wdata[9]\, sample_f0_wdata_10 => 
        \sample_f0_wdata[10]\, sample_f0_wdata_11 => 
        \sample_f0_wdata[11]\, sample_f0_wdata_12 => 
        \sample_f0_wdata[12]\, sample_f0_wdata_13 => 
        \sample_f0_wdata[13]\, sample_f0_wdata_14 => 
        \sample_f0_wdata[14]\, sample_f0_wdata_15 => 
        \sample_f0_wdata[15]\, sample_f0_wdata_48 => 
        \sample_f0_wdata[48]\, sample_f0_wdata_49 => 
        \sample_f0_wdata[49]\, sample_f0_wdata_50 => 
        \sample_f0_wdata[50]\, sample_f0_wdata_51 => 
        \sample_f0_wdata[51]\, sample_f0_wdata_52 => 
        \sample_f0_wdata[52]\, sample_f0_wdata_53 => 
        \sample_f0_wdata[53]\, sample_f0_wdata_54 => 
        \sample_f0_wdata[54]\, sample_f0_wdata_55 => 
        \sample_f0_wdata[55]\, sample_f0_wdata_56 => 
        \sample_f0_wdata[56]\, sample_f0_wdata_57 => 
        \sample_f0_wdata[57]\, sample_f0_wdata_58 => 
        \sample_f0_wdata[58]\, sample_f0_wdata_59 => 
        \sample_f0_wdata[59]\, sample_f0_wdata_60 => 
        \sample_f0_wdata[60]\, sample_f0_wdata_61 => 
        \sample_f0_wdata[61]\, sample_f0_wdata_62 => 
        \sample_f0_wdata[62]\, sample_f0_wdata_63 => 
        \sample_f0_wdata[63]\, sample_f0_wdata_64 => 
        \sample_f0_wdata[64]\, sample_f0_wdata_65 => 
        \sample_f0_wdata[65]\, sample_f0_wdata_66 => 
        \sample_f0_wdata[66]\, sample_f0_wdata_67 => 
        \sample_f0_wdata[67]\, sample_f0_wdata_68 => 
        \sample_f0_wdata[68]\, sample_f0_wdata_69 => 
        \sample_f0_wdata[69]\, sample_f0_wdata_70 => 
        \sample_f0_wdata[70]\, sample_f0_wdata_71 => 
        \sample_f0_wdata[71]\, sample_f0_wdata_72 => 
        \sample_f0_wdata[72]\, sample_f0_wdata_73 => 
        \sample_f0_wdata[73]\, sample_f0_wdata_74 => 
        \sample_f0_wdata[74]\, sample_f0_wdata_75 => 
        \sample_f0_wdata[75]\, sample_f0_wdata_76 => 
        \sample_f0_wdata[76]\, sample_f0_wdata_77 => 
        \sample_f0_wdata[77]\, sample_f0_wdata_78 => 
        \sample_f0_wdata[78]\, sample_f0_wdata_79 => 
        \sample_f0_wdata[79]\, sample_f0_wdata_80 => 
        \sample_f0_wdata[80]\, sample_f0_wdata_81 => 
        \sample_f0_wdata[81]\, sample_f0_wdata_82 => 
        \sample_f0_wdata[82]\, sample_f0_wdata_83 => 
        \sample_f0_wdata[83]\, sample_f0_wdata_84 => 
        \sample_f0_wdata[84]\, sample_f0_wdata_85 => 
        \sample_f0_wdata[85]\, sample_f0_wdata_86 => 
        \sample_f0_wdata[86]\, sample_f0_wdata_87 => 
        \sample_f0_wdata[87]\, sample_f0_wdata_88 => 
        \sample_f0_wdata[88]\, sample_f0_wdata_89 => 
        \sample_f0_wdata[89]\, sample_f0_wdata_90 => 
        \sample_f0_wdata[90]\, sample_f0_wdata_91 => 
        \sample_f0_wdata[91]\, sample_f0_wdata_92 => 
        \sample_f0_wdata[92]\, sample_f0_wdata_93 => 
        \sample_f0_wdata[93]\, sample_f0_wdata_94 => 
        \sample_f0_wdata[94]\, sample_f0_wdata_95 => 
        \sample_f0_wdata[95]\, delta_f2_f1(9) => delta_f2_f1(9), 
        delta_f2_f1(8) => delta_f2_f1(8), delta_f2_f1(7) => 
        delta_f2_f1(7), delta_f2_f1(6) => delta_f2_f1(6), 
        delta_f2_f1(5) => delta_f2_f1(5), delta_f2_f1(4) => 
        delta_f2_f1(4), delta_f2_f1(3) => delta_f2_f1(3), 
        delta_f2_f1(2) => delta_f2_f1(2), delta_f2_f1(1) => 
        delta_f2_f1(1), delta_f2_f1(0) => delta_f2_f1(0), 
        delta_snapshot(15) => delta_snapshot(15), 
        delta_snapshot(14) => delta_snapshot(14), 
        delta_snapshot(13) => delta_snapshot(13), 
        delta_snapshot(12) => delta_snapshot(12), 
        delta_snapshot(11) => delta_snapshot(11), 
        delta_snapshot(10) => delta_snapshot(10), 
        delta_snapshot(9) => delta_snapshot(9), delta_snapshot(8)
         => delta_snapshot(8), delta_snapshot(7) => 
        delta_snapshot(7), delta_snapshot(6) => delta_snapshot(6), 
        delta_snapshot(5) => delta_snapshot(5), delta_snapshot(4)
         => delta_snapshot(4), delta_snapshot(3) => 
        delta_snapshot(3), delta_snapshot(2) => delta_snapshot(2), 
        delta_snapshot(1) => delta_snapshot(1), delta_snapshot(0)
         => delta_snapshot(0), delta_f2_f0(9) => delta_f2_f0(9), 
        delta_f2_f0(8) => delta_f2_f0(8), delta_f2_f0(7) => 
        delta_f2_f0(7), delta_f2_f0(6) => delta_f2_f0(6), 
        delta_f2_f0(5) => delta_f2_f0(5), delta_f2_f0(4) => 
        delta_f2_f0(4), delta_f2_f0(3) => delta_f2_f0(3), 
        delta_f2_f0(2) => delta_f2_f0(2), delta_f2_f0(1) => 
        delta_f2_f0(1), delta_f2_f0(0) => delta_f2_f0(0), 
        nb_snapshot_param(10) => nb_snapshot_param(10), 
        nb_snapshot_param(9) => nb_snapshot_param(9), 
        nb_snapshot_param(8) => nb_snapshot_param(8), 
        nb_snapshot_param(7) => nb_snapshot_param(7), 
        nb_snapshot_param(6) => nb_snapshot_param(6), 
        nb_snapshot_param(5) => nb_snapshot_param(5), 
        nb_snapshot_param(4) => nb_snapshot_param(4), 
        nb_snapshot_param(3) => nb_snapshot_param(3), 
        nb_snapshot_param(2) => nb_snapshot_param(2), 
        nb_snapshot_param(1) => nb_snapshot_param(1), 
        nb_snapshot_param(0) => nb_snapshot_param(0), hwrite_c
         => hwrite_c, IdlePhase_RNI03G71 => IdlePhase_RNI03G71, 
        N_43 => N_43, lpp_waveform_GND => 
        lpp_top_lfr_wf_picker_ip_GND, lpp_waveform_VCC => 
        lpp_top_lfr_wf_picker_ip_VCC, sample_f3_val => 
        sample_f3_val, enable_f3 => enable_f3, burst_f2 => 
        burst_f2, enable_f2 => enable_f2, sample_f1_val_0 => 
        sample_f1_val_0, burst_f1 => burst_f1, enable_f1 => 
        enable_f1, data_shaping_R1_0 => data_shaping_R1_0, 
        data_shaping_R1 => data_shaping_R1, burst_f0 => burst_f0, 
        data_shaping_R0_0 => data_shaping_R0_0, data_shaping_R0
         => data_shaping_R0, enable_f0 => enable_f0, 
        coarse_time_0_c => coarse_time_0_c, sample_f2_val => 
        sample_f2_val, sample_f0_val_0 => sample_f0_val_0, HCLK_c
         => HCLK_c, HRESETn_c => HRESETn_c);
    
    Downsampling_f0 : Downsampling_8_16_4
      port map(sample_f0_0 => \sample_f0[48]\, sample_f0_1 => 
        \sample_f0[49]\, sample_f0_2 => \sample_f0[50]\, 
        sample_f0_3 => \sample_f0[51]\, sample_f0_4 => 
        \sample_f0[52]\, sample_f0_5 => \sample_f0[53]\, 
        sample_f0_6 => \sample_f0[54]\, sample_f0_7 => 
        \sample_f0[55]\, sample_f0_8 => \sample_f0[56]\, 
        sample_f0_9 => \sample_f0[57]\, sample_f0_10 => 
        \sample_f0[58]\, sample_f0_11 => \sample_f0[59]\, 
        sample_f0_12 => \sample_f0[60]\, sample_f0_13 => 
        \sample_f0[61]\, sample_f0_14 => \sample_f0[62]\, 
        sample_f0_15 => \sample_f0[63]\, sample_f0_32 => 
        \sample_f0[80]\, sample_f0_33 => \sample_f0[81]\, 
        sample_f0_34 => \sample_f0[82]\, sample_f0_35 => 
        \sample_f0[83]\, sample_f0_36 => \sample_f0[84]\, 
        sample_f0_37 => \sample_f0[85]\, sample_f0_38 => 
        \sample_f0[86]\, sample_f0_39 => \sample_f0[87]\, 
        sample_f0_40 => \sample_f0[88]\, sample_f0_41 => 
        \sample_f0[89]\, sample_f0_42 => \sample_f0[90]\, 
        sample_f0_43 => \sample_f0[91]\, sample_f0_44 => 
        \sample_f0[92]\, sample_f0_45 => \sample_f0[93]\, 
        sample_f0_46 => \sample_f0[94]\, sample_f0_47 => 
        \sample_f0[95]\, sample_f0_48 => \sample_f0[96]\, 
        sample_f0_49 => \sample_f0[97]\, sample_f0_50 => 
        \sample_f0[98]\, sample_f0_51 => \sample_f0[99]\, 
        sample_f0_52 => \sample_f0[100]\, sample_f0_53 => 
        \sample_f0[101]\, sample_f0_54 => \sample_f0[102]\, 
        sample_f0_55 => \sample_f0[103]\, sample_f0_56 => 
        \sample_f0[104]\, sample_f0_57 => \sample_f0[105]\, 
        sample_f0_58 => \sample_f0[106]\, sample_f0_59 => 
        \sample_f0[107]\, sample_f0_60 => \sample_f0[108]\, 
        sample_f0_61 => \sample_f0[109]\, sample_f0_62 => 
        \sample_f0[110]\, sample_f0_63 => \sample_f0[111]\, 
        sample_data_shaping_out_0 => \sample_data_shaping_out[2]\, 
        sample_data_shaping_out_1 => \sample_data_shaping_out[3]\, 
        sample_data_shaping_out_2 => \sample_data_shaping_out[4]\, 
        sample_data_shaping_out_3 => \sample_data_shaping_out[5]\, 
        sample_data_shaping_out_4 => \sample_data_shaping_out[6]\, 
        sample_data_shaping_out_5 => \sample_data_shaping_out[7]\, 
        sample_data_shaping_out_6 => \sample_data_shaping_out[8]\, 
        sample_data_shaping_out_7 => \sample_data_shaping_out[9]\, 
        sample_data_shaping_out_8 => 
        \sample_data_shaping_out[10]\, sample_data_shaping_out_9
         => \sample_data_shaping_out[11]\, 
        sample_data_shaping_out_10 => 
        \sample_data_shaping_out[12]\, sample_data_shaping_out_11
         => \sample_data_shaping_out[13]\, 
        sample_data_shaping_out_12 => 
        \sample_data_shaping_out[14]\, sample_data_shaping_out_13
         => \sample_data_shaping_out[15]\, 
        sample_data_shaping_out_14 => 
        \sample_data_shaping_out[16]\, sample_data_shaping_out_15
         => \sample_data_shaping_out[17]\, 
        sample_data_shaping_out_18 => 
        \sample_data_shaping_out[20]\, sample_data_shaping_out_19
         => \sample_data_shaping_out[21]\, 
        sample_data_shaping_out_20 => 
        \sample_data_shaping_out[22]\, sample_data_shaping_out_21
         => \sample_data_shaping_out[23]\, 
        sample_data_shaping_out_22 => 
        \sample_data_shaping_out[24]\, sample_data_shaping_out_23
         => \sample_data_shaping_out[25]\, 
        sample_data_shaping_out_24 => 
        \sample_data_shaping_out[26]\, sample_data_shaping_out_25
         => \sample_data_shaping_out[27]\, 
        sample_data_shaping_out_26 => 
        \sample_data_shaping_out[28]\, sample_data_shaping_out_27
         => \sample_data_shaping_out[29]\, 
        sample_data_shaping_out_28 => 
        \sample_data_shaping_out[30]\, sample_data_shaping_out_29
         => \sample_data_shaping_out[31]\, 
        sample_data_shaping_out_30 => 
        \sample_data_shaping_out[32]\, sample_data_shaping_out_31
         => \sample_data_shaping_out[33]\, 
        sample_data_shaping_out_32 => 
        \sample_data_shaping_out[34]\, sample_data_shaping_out_33
         => \sample_data_shaping_out[35]\, 
        sample_data_shaping_out_36 => 
        \sample_data_shaping_out[38]\, sample_data_shaping_out_37
         => \sample_data_shaping_out[39]\, 
        sample_data_shaping_out_38 => 
        \sample_data_shaping_out[40]\, sample_data_shaping_out_39
         => \sample_data_shaping_out[41]\, 
        sample_data_shaping_out_40 => 
        \sample_data_shaping_out[42]\, sample_data_shaping_out_41
         => \sample_data_shaping_out[43]\, 
        sample_data_shaping_out_42 => 
        \sample_data_shaping_out[44]\, sample_data_shaping_out_43
         => \sample_data_shaping_out[45]\, 
        sample_data_shaping_out_44 => 
        \sample_data_shaping_out[46]\, sample_data_shaping_out_45
         => \sample_data_shaping_out[47]\, 
        sample_data_shaping_out_46 => 
        \sample_data_shaping_out[48]\, sample_data_shaping_out_47
         => \sample_data_shaping_out[49]\, 
        sample_data_shaping_out_48 => 
        \sample_data_shaping_out[50]\, sample_data_shaping_out_49
         => \sample_data_shaping_out[51]\, 
        sample_data_shaping_out_50 => 
        \sample_data_shaping_out[52]\, sample_data_shaping_out_51
         => \sample_data_shaping_out[53]\, 
        sample_data_shaping_out_54 => 
        \sample_data_shaping_out[56]\, sample_data_shaping_out_55
         => \sample_data_shaping_out[57]\, 
        sample_data_shaping_out_56 => 
        \sample_data_shaping_out[58]\, sample_data_shaping_out_57
         => \sample_data_shaping_out[59]\, 
        sample_data_shaping_out_58 => 
        \sample_data_shaping_out[60]\, sample_data_shaping_out_59
         => \sample_data_shaping_out[61]\, 
        sample_data_shaping_out_60 => 
        \sample_data_shaping_out[62]\, sample_data_shaping_out_61
         => \sample_data_shaping_out[63]\, 
        sample_data_shaping_out_62 => 
        \sample_data_shaping_out[64]\, sample_data_shaping_out_63
         => \sample_data_shaping_out[65]\, 
        sample_data_shaping_out_64 => 
        \sample_data_shaping_out[66]\, sample_data_shaping_out_65
         => \sample_data_shaping_out[67]\, 
        sample_data_shaping_out_66 => 
        \sample_data_shaping_out[68]\, sample_data_shaping_out_67
         => \sample_data_shaping_out[69]\, 
        sample_data_shaping_out_68 => 
        \sample_data_shaping_out[70]\, sample_data_shaping_out_69
         => \sample_data_shaping_out[71]\, 
        sample_data_shaping_out_90 => 
        \sample_data_shaping_out[92]\, sample_data_shaping_out_91
         => \sample_data_shaping_out[93]\, 
        sample_data_shaping_out_92 => 
        \sample_data_shaping_out[94]\, sample_data_shaping_out_93
         => \sample_data_shaping_out[95]\, 
        sample_data_shaping_out_94 => 
        \sample_data_shaping_out[96]\, sample_data_shaping_out_95
         => \sample_data_shaping_out[97]\, 
        sample_data_shaping_out_96 => 
        \sample_data_shaping_out[98]\, sample_data_shaping_out_97
         => \sample_data_shaping_out[99]\, 
        sample_data_shaping_out_98 => 
        \sample_data_shaping_out[100]\, 
        sample_data_shaping_out_99 => 
        \sample_data_shaping_out[101]\, 
        sample_data_shaping_out_100 => 
        \sample_data_shaping_out[102]\, 
        sample_data_shaping_out_101 => 
        \sample_data_shaping_out[103]\, 
        sample_data_shaping_out_102 => 
        \sample_data_shaping_out[104]\, 
        sample_data_shaping_out_103 => 
        \sample_data_shaping_out[105]\, 
        sample_data_shaping_out_104 => 
        \sample_data_shaping_out[106]\, 
        sample_data_shaping_out_105 => 
        \sample_data_shaping_out[107]\, 
        sample_data_shaping_out_108 => 
        \sample_data_shaping_out[110]\, 
        sample_data_shaping_out_109 => 
        \sample_data_shaping_out[111]\, 
        sample_data_shaping_out_110 => 
        \sample_data_shaping_out[112]\, 
        sample_data_shaping_out_111 => 
        \sample_data_shaping_out[113]\, 
        sample_data_shaping_out_112 => 
        \sample_data_shaping_out[114]\, 
        sample_data_shaping_out_113 => 
        \sample_data_shaping_out[115]\, 
        sample_data_shaping_out_114 => 
        \sample_data_shaping_out[116]\, 
        sample_data_shaping_out_115 => 
        \sample_data_shaping_out[117]\, 
        sample_data_shaping_out_116 => 
        \sample_data_shaping_out[118]\, 
        sample_data_shaping_out_117 => 
        \sample_data_shaping_out[119]\, 
        sample_data_shaping_out_118 => 
        \sample_data_shaping_out[120]\, 
        sample_data_shaping_out_119 => 
        \sample_data_shaping_out[121]\, 
        sample_data_shaping_out_120 => 
        \sample_data_shaping_out[122]\, 
        sample_data_shaping_out_121 => 
        \sample_data_shaping_out[123]\, 
        sample_data_shaping_out_122 => 
        \sample_data_shaping_out[124]\, 
        sample_data_shaping_out_123 => 
        \sample_data_shaping_out[125]\, 
        sample_data_shaping_out_126 => 
        \sample_data_shaping_out[128]\, 
        sample_data_shaping_out_127 => 
        \sample_data_shaping_out[129]\, 
        sample_data_shaping_out_128 => 
        \sample_data_shaping_out[130]\, 
        sample_data_shaping_out_129 => 
        \sample_data_shaping_out[131]\, 
        sample_data_shaping_out_130 => 
        \sample_data_shaping_out[132]\, 
        sample_data_shaping_out_131 => 
        \sample_data_shaping_out[133]\, 
        sample_data_shaping_out_132 => 
        \sample_data_shaping_out[134]\, 
        sample_data_shaping_out_133 => 
        \sample_data_shaping_out[135]\, 
        sample_data_shaping_out_134 => 
        \sample_data_shaping_out[136]\, 
        sample_data_shaping_out_135 => 
        \sample_data_shaping_out[137]\, 
        sample_data_shaping_out_136 => 
        \sample_data_shaping_out[138]\, 
        sample_data_shaping_out_137 => 
        \sample_data_shaping_out[139]\, 
        sample_data_shaping_out_138 => 
        \sample_data_shaping_out[140]\, 
        sample_data_shaping_out_139 => 
        \sample_data_shaping_out[141]\, 
        sample_data_shaping_out_140 => 
        \sample_data_shaping_out[142]\, 
        sample_data_shaping_out_141 => 
        \sample_data_shaping_out[143]\, sample_f0_wdata_95 => 
        \sample_f0_wdata[95]\, sample_f0_wdata_94 => 
        \sample_f0_wdata[94]\, sample_f0_wdata_93 => 
        \sample_f0_wdata[93]\, sample_f0_wdata_92 => 
        \sample_f0_wdata[92]\, sample_f0_wdata_91 => 
        \sample_f0_wdata[91]\, sample_f0_wdata_90 => 
        \sample_f0_wdata[90]\, sample_f0_wdata_89 => 
        \sample_f0_wdata[89]\, sample_f0_wdata_88 => 
        \sample_f0_wdata[88]\, sample_f0_wdata_87 => 
        \sample_f0_wdata[87]\, sample_f0_wdata_86 => 
        \sample_f0_wdata[86]\, sample_f0_wdata_85 => 
        \sample_f0_wdata[85]\, sample_f0_wdata_84 => 
        \sample_f0_wdata[84]\, sample_f0_wdata_83 => 
        \sample_f0_wdata[83]\, sample_f0_wdata_82 => 
        \sample_f0_wdata[82]\, sample_f0_wdata_81 => 
        \sample_f0_wdata[81]\, sample_f0_wdata_80 => 
        \sample_f0_wdata[80]\, sample_f0_wdata_79 => 
        \sample_f0_wdata[79]\, sample_f0_wdata_78 => 
        \sample_f0_wdata[78]\, sample_f0_wdata_77 => 
        \sample_f0_wdata[77]\, sample_f0_wdata_76 => 
        \sample_f0_wdata[76]\, sample_f0_wdata_75 => 
        \sample_f0_wdata[75]\, sample_f0_wdata_74 => 
        \sample_f0_wdata[74]\, sample_f0_wdata_73 => 
        \sample_f0_wdata[73]\, sample_f0_wdata_72 => 
        \sample_f0_wdata[72]\, sample_f0_wdata_71 => 
        \sample_f0_wdata[71]\, sample_f0_wdata_70 => 
        \sample_f0_wdata[70]\, sample_f0_wdata_69 => 
        \sample_f0_wdata[69]\, sample_f0_wdata_68 => 
        \sample_f0_wdata[68]\, sample_f0_wdata_67 => 
        \sample_f0_wdata[67]\, sample_f0_wdata_66 => 
        \sample_f0_wdata[66]\, sample_f0_wdata_65 => 
        \sample_f0_wdata[65]\, sample_f0_wdata_64 => 
        \sample_f0_wdata[64]\, sample_f0_wdata_63 => 
        \sample_f0_wdata[63]\, sample_f0_wdata_62 => 
        \sample_f0_wdata[62]\, sample_f0_wdata_61 => 
        \sample_f0_wdata[61]\, sample_f0_wdata_60 => 
        \sample_f0_wdata[60]\, sample_f0_wdata_59 => 
        \sample_f0_wdata[59]\, sample_f0_wdata_58 => 
        \sample_f0_wdata[58]\, sample_f0_wdata_57 => 
        \sample_f0_wdata[57]\, sample_f0_wdata_56 => 
        \sample_f0_wdata[56]\, sample_f0_wdata_55 => 
        \sample_f0_wdata[55]\, sample_f0_wdata_54 => 
        \sample_f0_wdata[54]\, sample_f0_wdata_53 => 
        \sample_f0_wdata[53]\, sample_f0_wdata_52 => 
        \sample_f0_wdata[52]\, sample_f0_wdata_51 => 
        \sample_f0_wdata[51]\, sample_f0_wdata_50 => 
        \sample_f0_wdata[50]\, sample_f0_wdata_49 => 
        \sample_f0_wdata[49]\, sample_f0_wdata_48 => 
        \sample_f0_wdata[48]\, sample_f0_wdata_15 => 
        \sample_f0_wdata[15]\, sample_f0_wdata_14 => 
        \sample_f0_wdata[14]\, sample_f0_wdata_13 => 
        \sample_f0_wdata[13]\, sample_f0_wdata_12 => 
        \sample_f0_wdata[12]\, sample_f0_wdata_11 => 
        \sample_f0_wdata[11]\, sample_f0_wdata_10 => 
        \sample_f0_wdata[10]\, sample_f0_wdata_9 => 
        \sample_f0_wdata[9]\, sample_f0_wdata_8 => 
        \sample_f0_wdata[8]\, sample_f0_wdata_7 => 
        \sample_f0_wdata[7]\, sample_f0_wdata_6 => 
        \sample_f0_wdata[6]\, sample_f0_wdata_5 => 
        \sample_f0_wdata[5]\, sample_f0_wdata_4 => 
        \sample_f0_wdata[4]\, sample_f0_wdata_3 => 
        \sample_f0_wdata[3]\, sample_f0_wdata_2 => 
        \sample_f0_wdata[2]\, sample_f0_wdata_1 => 
        \sample_f0_wdata[1]\, sample_f0_wdata_0 => 
        \sample_f0_wdata[0]\, sample_data_shaping_out_val => 
        \sample_data_shaping_out_val\, sample_f0_val => 
        sample_f0_val, sample_data_shaping_out_val_0 => 
        \sample_data_shaping_out_val_0\, sample_f0_val_0 => 
        sample_f0_val_0, HRESETn_c => HRESETn_c, HCLK_c => HCLK_c, 
        sample_f0_val_1 => sample_f0_val_1);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[51]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[51]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[51]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[141]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[141]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[141]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I95_Y_0 : 
        AX1D
      port map(A => I92_un1_Y, B => N182_0, C => N183, Y => 
        \sample_data_shaping_f1_f0_s[2]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I37_Y : 
        XA1A
      port map(A => \sample_filter_v2_out[115]\, B => 
        \sample_filter_v2_out[133]\, C => N197, Y => N216);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out_RNO[106]\ : 
        MX2
      port map(A => \sample_filter_v2_out[106]\, B => 
        \sample_data_shaping_f2_f1_s[1]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_41[106]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I49_Y : 
        AO1B
      port map(A => N264_0, B => N216_0, C => 
        SUB_16x16_medium_area_I49_Y_0, Y => N244);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I57_Y_0 : 
        AO18
      port map(A => N206_0, B => \sample_filter_v2_out[129]\, C
         => \sample_filter_v2_out[111]\, Y => 
        SUB_16x16_medium_area_I57_Y_0_0);
    
    sample_data_shaping_out_val : DFN1C0
      port map(D => sample_filter_v2_out_val, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out_val\);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out_RNO[125]\ : 
        AX1C
      port map(A => \sample_filter_v2_out[143]\, B => 
        data_shaping_SP0, C => \sample_filter_v2_out[125]\, Y => 
        \sample_data_shaping_out_13[125]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I103_Y_0 : 
        AX1D
      port map(A => I88_un1_Y, B => N198, C => N199, Y => 
        \sample_data_shaping_f2_f1_s[10]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I23_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[118]\, B => 
        \sample_filter_v2_out[136]\, Y => N194);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[106]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_41[106]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[106]\);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[118]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_181[118]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[118]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I99_Y_0 : 
        XOR3
      port map(A => \sample_filter_v2_out[101]\, B => 
        \sample_filter_v2_out[119]\, C => N290_i, Y => 
        \sample_data_shaping_f2_f1_s[6]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[102]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_137[102]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[102]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I90_un1_Y : 
        OA1
      port map(A => I85_un1_Y, B => N274_0, C => N189, Y => 
        I90_un1_Y);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I46_Y : 
        OR2A
      port map(A => \sample_filter_v2_out[125]\, B => 
        \sample_filter_v2_out[107]\, Y => N225);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[4]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[4]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[4]\);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[125]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_13[125]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[125]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I99_Y_0 : 
        AX1D
      port map(A => I90_un1_Y, B => N190_0, C => N191, Y => 
        \sample_data_shaping_f1_f0_s[6]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I29_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[130]\, B => 
        \sample_filter_v2_out[112]\, Y => N205);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[6]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[6]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[6]\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[69]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[69]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[69]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[25]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[25]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[25]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[121]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_109[121]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[121]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I90_Y : 
        AO18
      port map(A => N280, B => \sample_filter_v2_out[120]\, C => 
        \sample_filter_v2_out[102]\, Y => N290_i);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[94]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_329[94]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[94]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I57_Y_1 : 
        OA1
      port map(A => N212_0, B => N254_0, C => 
        SUB_16x16_medium_area_I57_Y_0_0, Y => 
        SUB_16x16_medium_area_I57_Y_1_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I39_Y : 
        NOR2B
      port map(A => N195_0, B => N193, Y => N265_0);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[53]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[53]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[53]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I57_Y_0 : 
        AO18
      port map(A => N206, B => \sample_filter_v2_out[111]\, C => 
        \sample_filter_v2_out[93]\, Y => 
        SUB_16x16_medium_area_I57_Y_0);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out_RNO[124]\ : 
        MX2
      port map(A => \sample_filter_v2_out[124]\, B => 
        \sample_data_shaping_f1_f0_s[1]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_37[124]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I108_Y_0 : 
        XNOR3
      port map(A => \sample_filter_v2_out[110]\, B => 
        \sample_filter_v2_out[92]\, C => N240_0, Y => 
        \sample_data_shaping_f2_f1_s[15]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I94_Y_0 : 
        XOR2
      port map(A => N225, B => N181_0, Y => 
        \sample_data_shaping_f2_f1_s[1]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I29_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[112]\, B => 
        \sample_filter_v2_out[130]\, Y => N206_0);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[99]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_209[99]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[99]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I88_Y : 
        AO18
      port map(A => N270, B => \sample_filter_v2_out[134]\, C => 
        \sample_filter_v2_out[116]\, Y => N286_i);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[116]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_229[116]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[116]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I50_Y : 
        NOR2B
      port map(A => N265, B => N216, Y => N245_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I24_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[117]\, B => 
        \sample_filter_v2_out[99]\, Y => N195_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I18_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[141]\, B => 
        \sample_filter_v2_out[123]\, Y => N183);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out_RNO[119]\ : 
        MX2
      port map(A => \sample_filter_v2_out[119]\, B => 
        \sample_data_shaping_f1_f0_s[6]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_157[119]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[139]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[139]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[139]\);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[70]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[70]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[70]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I27_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[114]\, B => 
        \sample_filter_v2_out[96]\, Y => N201_0);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[8]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[8]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[8]\);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[112]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_325[112]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[112]\);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[98]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_233[98]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[98]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[128]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[128]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[128]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I56_Y_0 : 
        AO18
      port map(A => N190, B => \sample_filter_v2_out[119]\, C => 
        \sample_filter_v2_out[101]\, Y => 
        SUB_16x16_medium_area_I56_Y_0);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[134]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[134]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[134]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I25_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[116]\, B => 
        \sample_filter_v2_out[98]\, Y => N197_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I29_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[112]\, B => 
        \sample_filter_v2_out[94]\, Y => N205_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I64_Y : 
        AO1
      port map(A => N268, B => N245_0, C => N244_0, Y => N258);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I57_Y : 
        AO1B
      port map(A => SUB_16x16_medium_area_I57_un1_Y_0_0, B => 
        N268, C => SUB_16x16_medium_area_I57_Y_2_0, Y => N240);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[59]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[59]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[59]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I34_Y : 
        AO13
      port map(A => N202_0, B => \sample_filter_v2_out[95]\, C
         => \sample_filter_v2_out[113]\, Y => N254);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[10]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[10]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[10]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I96_Y_0 : 
        XOR2
      port map(A => N278, B => N185, Y => 
        \sample_data_shaping_f1_f0_s[3]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I21_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[120]\, B => 
        \sample_filter_v2_out[138]\, Y => N190_0);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[40]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[40]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[40]\);
    
    Downsampling_f1 : Downsampling_8_16_6
      port map(sample_f0_0 => \sample_f0[48]\, sample_f0_1 => 
        \sample_f0[49]\, sample_f0_2 => \sample_f0[50]\, 
        sample_f0_3 => \sample_f0[51]\, sample_f0_4 => 
        \sample_f0[52]\, sample_f0_5 => \sample_f0[53]\, 
        sample_f0_6 => \sample_f0[54]\, sample_f0_7 => 
        \sample_f0[55]\, sample_f0_8 => \sample_f0[56]\, 
        sample_f0_9 => \sample_f0[57]\, sample_f0_10 => 
        \sample_f0[58]\, sample_f0_11 => \sample_f0[59]\, 
        sample_f0_12 => \sample_f0[60]\, sample_f0_13 => 
        \sample_f0[61]\, sample_f0_14 => \sample_f0[62]\, 
        sample_f0_15 => \sample_f0[63]\, sample_f0_32 => 
        \sample_f0[80]\, sample_f0_33 => \sample_f0[81]\, 
        sample_f0_34 => \sample_f0[82]\, sample_f0_35 => 
        \sample_f0[83]\, sample_f0_36 => \sample_f0[84]\, 
        sample_f0_37 => \sample_f0[85]\, sample_f0_38 => 
        \sample_f0[86]\, sample_f0_39 => \sample_f0[87]\, 
        sample_f0_40 => \sample_f0[88]\, sample_f0_41 => 
        \sample_f0[89]\, sample_f0_42 => \sample_f0[90]\, 
        sample_f0_43 => \sample_f0[91]\, sample_f0_44 => 
        \sample_f0[92]\, sample_f0_45 => \sample_f0[93]\, 
        sample_f0_46 => \sample_f0[94]\, sample_f0_47 => 
        \sample_f0[95]\, sample_f0_48 => \sample_f0[96]\, 
        sample_f0_49 => \sample_f0[97]\, sample_f0_50 => 
        \sample_f0[98]\, sample_f0_51 => \sample_f0[99]\, 
        sample_f0_52 => \sample_f0[100]\, sample_f0_53 => 
        \sample_f0[101]\, sample_f0_54 => \sample_f0[102]\, 
        sample_f0_55 => \sample_f0[103]\, sample_f0_56 => 
        \sample_f0[104]\, sample_f0_57 => \sample_f0[105]\, 
        sample_f0_58 => \sample_f0[106]\, sample_f0_59 => 
        \sample_f0[107]\, sample_f0_60 => \sample_f0[108]\, 
        sample_f0_61 => \sample_f0[109]\, sample_f0_62 => 
        \sample_f0[110]\, sample_f0_63 => \sample_f0[111]\, 
        sample_f1_0 => \sample_f1[48]\, sample_f1_1 => 
        \sample_f1[49]\, sample_f1_2 => \sample_f1[50]\, 
        sample_f1_3 => \sample_f1[51]\, sample_f1_4 => 
        \sample_f1[52]\, sample_f1_5 => \sample_f1[53]\, 
        sample_f1_6 => \sample_f1[54]\, sample_f1_7 => 
        \sample_f1[55]\, sample_f1_8 => \sample_f1[56]\, 
        sample_f1_9 => \sample_f1[57]\, sample_f1_10 => 
        \sample_f1[58]\, sample_f1_11 => \sample_f1[59]\, 
        sample_f1_12 => \sample_f1[60]\, sample_f1_13 => 
        \sample_f1[61]\, sample_f1_14 => \sample_f1[62]\, 
        sample_f1_15 => \sample_f1[63]\, sample_f1_32 => 
        \sample_f1[80]\, sample_f1_33 => \sample_f1[81]\, 
        sample_f1_34 => \sample_f1[82]\, sample_f1_35 => 
        \sample_f1[83]\, sample_f1_36 => \sample_f1[84]\, 
        sample_f1_37 => \sample_f1[85]\, sample_f1_38 => 
        \sample_f1[86]\, sample_f1_39 => \sample_f1[87]\, 
        sample_f1_40 => \sample_f1[88]\, sample_f1_41 => 
        \sample_f1[89]\, sample_f1_42 => \sample_f1[90]\, 
        sample_f1_43 => \sample_f1[91]\, sample_f1_44 => 
        \sample_f1[92]\, sample_f1_45 => \sample_f1[93]\, 
        sample_f1_46 => \sample_f1[94]\, sample_f1_47 => 
        \sample_f1[95]\, sample_f1_48 => \sample_f1[96]\, 
        sample_f1_49 => \sample_f1[97]\, sample_f1_50 => 
        \sample_f1[98]\, sample_f1_51 => \sample_f1[99]\, 
        sample_f1_52 => \sample_f1[100]\, sample_f1_53 => 
        \sample_f1[101]\, sample_f1_54 => \sample_f1[102]\, 
        sample_f1_55 => \sample_f1[103]\, sample_f1_56 => 
        \sample_f1[104]\, sample_f1_57 => \sample_f1[105]\, 
        sample_f1_58 => \sample_f1[106]\, sample_f1_59 => 
        \sample_f1[107]\, sample_f1_60 => \sample_f1[108]\, 
        sample_f1_61 => \sample_f1[109]\, sample_f1_62 => 
        \sample_f1[110]\, sample_f1_63 => \sample_f1[111]\, 
        sample_f0_wdata_95 => \sample_f0_wdata[95]\, 
        sample_f0_wdata_94 => \sample_f0_wdata[94]\, 
        sample_f0_wdata_93 => \sample_f0_wdata[93]\, 
        sample_f0_wdata_92 => \sample_f0_wdata[92]\, 
        sample_f0_wdata_91 => \sample_f0_wdata[91]\, 
        sample_f0_wdata_90 => \sample_f0_wdata[90]\, 
        sample_f0_wdata_89 => \sample_f0_wdata[89]\, 
        sample_f0_wdata_88 => \sample_f0_wdata[88]\, 
        sample_f0_wdata_87 => \sample_f0_wdata[87]\, 
        sample_f0_wdata_86 => \sample_f0_wdata[86]\, 
        sample_f0_wdata_85 => \sample_f0_wdata[85]\, 
        sample_f0_wdata_84 => \sample_f0_wdata[84]\, 
        sample_f0_wdata_83 => \sample_f0_wdata[83]\, 
        sample_f0_wdata_82 => \sample_f0_wdata[82]\, 
        sample_f0_wdata_81 => \sample_f0_wdata[81]\, 
        sample_f0_wdata_80 => \sample_f0_wdata[80]\, 
        sample_f0_wdata_79 => \sample_f0_wdata[79]\, 
        sample_f0_wdata_78 => \sample_f0_wdata[78]\, 
        sample_f0_wdata_77 => \sample_f0_wdata[77]\, 
        sample_f0_wdata_76 => \sample_f0_wdata[76]\, 
        sample_f0_wdata_75 => \sample_f0_wdata[75]\, 
        sample_f0_wdata_74 => \sample_f0_wdata[74]\, 
        sample_f0_wdata_73 => \sample_f0_wdata[73]\, 
        sample_f0_wdata_72 => \sample_f0_wdata[72]\, 
        sample_f0_wdata_71 => \sample_f0_wdata[71]\, 
        sample_f0_wdata_70 => \sample_f0_wdata[70]\, 
        sample_f0_wdata_69 => \sample_f0_wdata[69]\, 
        sample_f0_wdata_68 => \sample_f0_wdata[68]\, 
        sample_f0_wdata_67 => \sample_f0_wdata[67]\, 
        sample_f0_wdata_66 => \sample_f0_wdata[66]\, 
        sample_f0_wdata_65 => \sample_f0_wdata[65]\, 
        sample_f0_wdata_64 => \sample_f0_wdata[64]\, 
        sample_f0_wdata_63 => \sample_f0_wdata[63]\, 
        sample_f0_wdata_62 => \sample_f0_wdata[62]\, 
        sample_f0_wdata_61 => \sample_f0_wdata[61]\, 
        sample_f0_wdata_60 => \sample_f0_wdata[60]\, 
        sample_f0_wdata_59 => \sample_f0_wdata[59]\, 
        sample_f0_wdata_58 => \sample_f0_wdata[58]\, 
        sample_f0_wdata_57 => \sample_f0_wdata[57]\, 
        sample_f0_wdata_56 => \sample_f0_wdata[56]\, 
        sample_f0_wdata_55 => \sample_f0_wdata[55]\, 
        sample_f0_wdata_54 => \sample_f0_wdata[54]\, 
        sample_f0_wdata_53 => \sample_f0_wdata[53]\, 
        sample_f0_wdata_52 => \sample_f0_wdata[52]\, 
        sample_f0_wdata_51 => \sample_f0_wdata[51]\, 
        sample_f0_wdata_50 => \sample_f0_wdata[50]\, 
        sample_f0_wdata_49 => \sample_f0_wdata[49]\, 
        sample_f0_wdata_48 => \sample_f0_wdata[48]\, 
        sample_f0_wdata_15 => \sample_f0_wdata[15]\, 
        sample_f0_wdata_14 => \sample_f0_wdata[14]\, 
        sample_f0_wdata_13 => \sample_f0_wdata[13]\, 
        sample_f0_wdata_12 => \sample_f0_wdata[12]\, 
        sample_f0_wdata_11 => \sample_f0_wdata[11]\, 
        sample_f0_wdata_10 => \sample_f0_wdata[10]\, 
        sample_f0_wdata_9 => \sample_f0_wdata[9]\, 
        sample_f0_wdata_8 => \sample_f0_wdata[8]\, 
        sample_f0_wdata_7 => \sample_f0_wdata[7]\, 
        sample_f0_wdata_6 => \sample_f0_wdata[6]\, 
        sample_f0_wdata_5 => \sample_f0_wdata[5]\, 
        sample_f0_wdata_4 => \sample_f0_wdata[4]\, 
        sample_f0_wdata_3 => \sample_f0_wdata[3]\, 
        sample_f0_wdata_2 => \sample_f0_wdata[2]\, 
        sample_f0_wdata_1 => \sample_f0_wdata[1]\, 
        sample_f0_wdata_0 => \sample_f0_wdata[0]\, 
        sample_f1_wdata_95 => \sample_f1_wdata[95]\, 
        sample_f1_wdata_94 => \sample_f1_wdata[94]\, 
        sample_f1_wdata_93 => \sample_f1_wdata[93]\, 
        sample_f1_wdata_92 => \sample_f1_wdata[92]\, 
        sample_f1_wdata_91 => \sample_f1_wdata[91]\, 
        sample_f1_wdata_90 => \sample_f1_wdata[90]\, 
        sample_f1_wdata_89 => \sample_f1_wdata[89]\, 
        sample_f1_wdata_88 => \sample_f1_wdata[88]\, 
        sample_f1_wdata_87 => \sample_f1_wdata[87]\, 
        sample_f1_wdata_86 => \sample_f1_wdata[86]\, 
        sample_f1_wdata_85 => \sample_f1_wdata[85]\, 
        sample_f1_wdata_84 => \sample_f1_wdata[84]\, 
        sample_f1_wdata_83 => \sample_f1_wdata[83]\, 
        sample_f1_wdata_82 => \sample_f1_wdata[82]\, 
        sample_f1_wdata_81 => \sample_f1_wdata[81]\, 
        sample_f1_wdata_80 => \sample_f1_wdata[80]\, 
        sample_f1_wdata_79 => \sample_f1_wdata[79]\, 
        sample_f1_wdata_78 => \sample_f1_wdata[78]\, 
        sample_f1_wdata_77 => \sample_f1_wdata[77]\, 
        sample_f1_wdata_76 => \sample_f1_wdata[76]\, 
        sample_f1_wdata_75 => \sample_f1_wdata[75]\, 
        sample_f1_wdata_74 => \sample_f1_wdata[74]\, 
        sample_f1_wdata_73 => \sample_f1_wdata[73]\, 
        sample_f1_wdata_72 => \sample_f1_wdata[72]\, 
        sample_f1_wdata_71 => \sample_f1_wdata[71]\, 
        sample_f1_wdata_70 => \sample_f1_wdata[70]\, 
        sample_f1_wdata_69 => \sample_f1_wdata[69]\, 
        sample_f1_wdata_68 => \sample_f1_wdata[68]\, 
        sample_f1_wdata_67 => \sample_f1_wdata[67]\, 
        sample_f1_wdata_66 => \sample_f1_wdata[66]\, 
        sample_f1_wdata_65 => \sample_f1_wdata[65]\, 
        sample_f1_wdata_64 => \sample_f1_wdata[64]\, 
        sample_f1_wdata_63 => \sample_f1_wdata[63]\, 
        sample_f1_wdata_62 => \sample_f1_wdata[62]\, 
        sample_f1_wdata_61 => \sample_f1_wdata[61]\, 
        sample_f1_wdata_60 => \sample_f1_wdata[60]\, 
        sample_f1_wdata_59 => \sample_f1_wdata[59]\, 
        sample_f1_wdata_58 => \sample_f1_wdata[58]\, 
        sample_f1_wdata_57 => \sample_f1_wdata[57]\, 
        sample_f1_wdata_56 => \sample_f1_wdata[56]\, 
        sample_f1_wdata_55 => \sample_f1_wdata[55]\, 
        sample_f1_wdata_54 => \sample_f1_wdata[54]\, 
        sample_f1_wdata_53 => \sample_f1_wdata[53]\, 
        sample_f1_wdata_52 => \sample_f1_wdata[52]\, 
        sample_f1_wdata_51 => \sample_f1_wdata[51]\, 
        sample_f1_wdata_50 => \sample_f1_wdata[50]\, 
        sample_f1_wdata_49 => \sample_f1_wdata[49]\, 
        sample_f1_wdata_48 => \sample_f1_wdata[48]\, 
        sample_f1_wdata_15 => \sample_f1_wdata[15]\, 
        sample_f1_wdata_14 => \sample_f1_wdata[14]\, 
        sample_f1_wdata_13 => \sample_f1_wdata[13]\, 
        sample_f1_wdata_12 => \sample_f1_wdata[12]\, 
        sample_f1_wdata_11 => \sample_f1_wdata[11]\, 
        sample_f1_wdata_10 => \sample_f1_wdata[10]\, 
        sample_f1_wdata_9 => \sample_f1_wdata[9]\, 
        sample_f1_wdata_8 => \sample_f1_wdata[8]\, 
        sample_f1_wdata_7 => \sample_f1_wdata[7]\, 
        sample_f1_wdata_6 => \sample_f1_wdata[6]\, 
        sample_f1_wdata_5 => \sample_f1_wdata[5]\, 
        sample_f1_wdata_4 => \sample_f1_wdata[4]\, 
        sample_f1_wdata_3 => \sample_f1_wdata[3]\, 
        sample_f1_wdata_2 => \sample_f1_wdata[2]\, 
        sample_f1_wdata_1 => \sample_f1_wdata[1]\, 
        sample_f1_wdata_0 => \sample_f1_wdata[0]\, 
        sample_f0_val_1 => sample_f0_val_1, sample_f1_val => 
        sample_f1_val, sample_f0_val_0 => sample_f0_val_0, 
        sample_out_0_sqmuxa_1 => sample_out_0_sqmuxa_1, HRESETn_c
         => HRESETn_c, HCLK_c => HCLK_c, sample_f1_val_0 => 
        sample_f1_val_0);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out_RNO[100]\ : 
        MX2
      port map(A => \sample_filter_v2_out[100]\, B => 
        \sample_data_shaping_f2_f1_s[7]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_185[100]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I49_Y : 
        AO1B
      port map(A => N264, B => N216, C => 
        SUB_16x16_medium_area_I49_Y_0_0, Y => N244_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I23_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[118]\, B => 
        \sample_filter_v2_out[100]\, Y => N193);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I41_Y : 
        XA1A
      port map(A => \sample_filter_v2_out[101]\, B => 
        \sample_filter_v2_out[119]\, C => N189_0, Y => N220);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I57_Y : 
        AO1B
      port map(A => SUB_16x16_medium_area_I57_un1_Y_0, B => 
        N268_0, C => SUB_16x16_medium_area_I57_Y_2, Y => N240_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I17_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[142]\, B => 
        \sample_filter_v2_out[124]\, Y => N181);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out_RNO[98]\ : 
        MX2
      port map(A => \sample_filter_v2_out[98]\, B => 
        \sample_data_shaping_f2_f1_s[9]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_233[98]\);
    
    sample_data_shaping_out_val_0 : DFN1C0
      port map(D => sample_filter_v2_out_val, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out_val_0\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I38_Y : 
        AO13
      port map(A => N194, B => \sample_filter_v2_out[117]\, C => 
        \sample_filter_v2_out[135]\, Y => N264);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[41]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[41]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[41]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[140]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[140]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[140]\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out_RNO[105]\ : 
        MX2
      port map(A => \sample_filter_v2_out[105]\, B => 
        \sample_data_shaping_f2_f1_s[2]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_65[105]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I57_Y_1 : 
        AOI1B
      port map(A => N254, B => N212, C => 
        SUB_16x16_medium_area_I57_Y_0, Y => 
        SUB_16x16_medium_area_I57_Y_1);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out_RNO[102]\ : 
        MX2
      port map(A => \sample_filter_v2_out[102]\, B => 
        \sample_data_shaping_f2_f1_s[5]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_137[102]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I57_Y_2 : 
        AOI1B
      port map(A => N244_0, B => N229_0, C => 
        SUB_16x16_medium_area_I57_Y_1_0, Y => 
        SUB_16x16_medium_area_I57_Y_2_0);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[39]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[39]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[39]\);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[130]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[130]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[130]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I97_Y_0 : 
        AX1D
      port map(A => SUB_16x16_medium_area_I91_un1_Y_0, B => 
        N186_0, C => N187_0, Y => 
        \sample_data_shaping_f2_f1_s[4]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I21_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[120]\, B => 
        \sample_filter_v2_out[102]\, Y => N189_0);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[63]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[63]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[63]\);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[101]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_161[101]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[101]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I106_Y_0 : 
        XOR2
      port map(A => N260, B => N205, Y => 
        \sample_data_shaping_f1_f0_s[13]\);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[45]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[45]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[45]\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[123]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_61[123]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[123]\);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[24]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[24]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[24]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out_RNO[122]\ : 
        MX2
      port map(A => \sample_filter_v2_out[122]\, B => 
        \sample_data_shaping_f1_f0_s[3]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_85[122]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[115]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_253[115]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[115]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[43]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[43]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[43]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I78_un1_Y : 
        NOR2B
      port map(A => N268_0, B => N265_0, Y => I78_un1_Y);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[60]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[60]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[60]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I42_Y : 
        AO13
      port map(A => N186, B => \sample_filter_v2_out[121]\, C => 
        \sample_filter_v2_out[139]\, Y => N274_0);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[64]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[64]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[64]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[133]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[133]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[133]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I57_Y_2 : 
        AOI1B
      port map(A => N244, B => N229, C => 
        SUB_16x16_medium_area_I57_Y_1, Y => 
        SUB_16x16_medium_area_I57_Y_2);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out_RNO[121]\ : 
        MX2
      port map(A => \sample_filter_v2_out[121]\, B => 
        \sample_data_shaping_f1_f0_s[4]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_109[121]\);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[142]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[142]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[142]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I96_Y_0 : 
        XNOR3
      port map(A => \sample_filter_v2_out[104]\, B => 
        \sample_filter_v2_out[122]\, C => N278_0, Y => 
        \sample_data_shaping_f2_f1_s[3]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I53_un1_Y : 
        OR3C
      port map(A => N225_0, B => N183, C => N181, Y => I53_un1_Y);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[14]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[14]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[14]\);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out_RNO[99]\ : 
        MX2
      port map(A => \sample_filter_v2_out[99]\, B => 
        \sample_data_shaping_f2_f1_s[8]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_209[99]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I101_Y_0 : 
        AX1D
      port map(A => SUB_16x16_medium_area_I89_un1_Y, B => N194_0, 
        C => N195_0, Y => \sample_data_shaping_f2_f1_s[8]\);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out_RNO[118]\ : 
        MX2
      port map(A => \sample_filter_v2_out[118]\, B => 
        \sample_data_shaping_f1_f0_s[7]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_181[118]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I103_Y_0 : 
        XOR3
      port map(A => \sample_filter_v2_out[115]\, B => 
        \sample_filter_v2_out[133]\, C => N286_i, Y => 
        \sample_data_shaping_f1_f0_s[10]\);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[93]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_353[93]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[93]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I92_un1_Y : 
        NOR2B
      port map(A => N225_0, B => N181, Y => I92_un1_Y);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out_RNO[117]\ : 
        MX2
      port map(A => \sample_filter_v2_out[117]\, B => 
        \sample_data_shaping_f1_f0_s[8]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_205[117]\);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out_RNO[112]\ : 
        MX2
      port map(A => \sample_filter_v2_out[112]\, B => 
        \sample_data_shaping_f1_f0_s[13]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_325[112]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I53_Y_0 : 
        AO18
      port map(A => N182, B => \sample_filter_v2_out[123]\, C => 
        \sample_filter_v2_out[105]\, Y => 
        SUB_16x16_medium_area_I53_Y_0);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[114]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_277[114]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[114]\);
    
    DIGITAL_acquisition : AD7688_drvr
      port map(sample_7(15) => \sample_7[15]\, sample_7(14) => 
        \sample_7[14]\, sample_7(13) => \sample_7[13]\, 
        sample_7(12) => \sample_7[12]\, sample_7(11) => 
        \sample_7[11]\, sample_7(10) => \sample_7[10]\, 
        sample_7(9) => \sample_7[9]\, sample_7(8) => 
        \sample_7[8]\, sample_7(7) => \sample_7[7]\, sample_7(6)
         => \sample_7[6]\, sample_7(5) => \sample_7[5]\, 
        sample_7(4) => \sample_7[4]\, sample_7(3) => 
        \sample_7[3]\, sample_7(2) => \sample_7[2]\, sample_7(1)
         => \sample_7[1]\, sample_7(0) => \sample_7[0]\, 
        sample_0(15) => \sample_0[15]\, sample_0(14) => 
        \sample_0[14]\, sample_0(13) => \sample_0[13]\, 
        sample_0(12) => \sample_0[12]\, sample_0(11) => 
        \sample_0[11]\, sample_0(10) => \sample_0[10]\, 
        sample_0(9) => \sample_0[9]\, sample_0(8) => 
        \sample_0[8]\, sample_0(7) => \sample_0[7]\, sample_0(6)
         => \sample_0[6]\, sample_0(5) => \sample_0[5]\, 
        sample_0(4) => \sample_0[4]\, sample_0(3) => 
        \sample_0[3]\, sample_0(2) => \sample_0[2]\, sample_0(1)
         => \sample_0[1]\, sample_0(0) => \sample_0[0]\, 
        sample_1(15) => \sample_1[15]\, sample_1(14) => 
        \sample_1[14]\, sample_1(13) => \sample_1[13]\, 
        sample_1(12) => \sample_1[12]\, sample_1(11) => 
        \sample_1[11]\, sample_1(10) => \sample_1[10]\, 
        sample_1(9) => \sample_1[9]\, sample_1(8) => 
        \sample_1[8]\, sample_1(7) => \sample_1[7]\, sample_1(6)
         => \sample_1[6]\, sample_1(5) => \sample_1[5]\, 
        sample_1(4) => \sample_1[4]\, sample_1(3) => 
        \sample_1[3]\, sample_1(2) => \sample_1[2]\, sample_1(1)
         => \sample_1[1]\, sample_1(0) => \sample_1[0]\, 
        sample_2(15) => \sample_2[15]\, sample_2(14) => 
        \sample_2[14]\, sample_2(13) => \sample_2[13]\, 
        sample_2(12) => \sample_2[12]\, sample_2(11) => 
        \sample_2[11]\, sample_2(10) => \sample_2[10]\, 
        sample_2(9) => \sample_2[9]\, sample_2(8) => 
        \sample_2[8]\, sample_2(7) => \sample_2[7]\, sample_2(6)
         => \sample_2[6]\, sample_2(5) => \sample_2[5]\, 
        sample_2(4) => \sample_2[4]\, sample_2(3) => 
        \sample_2[3]\, sample_2(2) => \sample_2[2]\, sample_2(1)
         => \sample_2[1]\, sample_2(0) => \sample_2[0]\, 
        sample_3(15) => \sample_3[15]\, sample_3(14) => 
        \sample_3[14]\, sample_3(13) => \sample_3[13]\, 
        sample_3(12) => \sample_3[12]\, sample_3(11) => 
        \sample_3[11]\, sample_3(10) => \sample_3[10]\, 
        sample_3(9) => \sample_3[9]\, sample_3(8) => 
        \sample_3[8]\, sample_3(7) => \sample_3[7]\, sample_3(6)
         => \sample_3[6]\, sample_3(5) => \sample_3[5]\, 
        sample_3(4) => \sample_3[4]\, sample_3(3) => 
        \sample_3[3]\, sample_3(2) => \sample_3[2]\, sample_3(1)
         => \sample_3[1]\, sample_3(0) => \sample_3[0]\, 
        sample_4(15) => \sample_4[15]\, sample_4(14) => 
        \sample_4[14]\, sample_4(13) => \sample_4[13]\, 
        sample_4(12) => \sample_4[12]\, sample_4(11) => 
        \sample_4[11]\, sample_4(10) => \sample_4[10]\, 
        sample_4(9) => \sample_4[9]\, sample_4(8) => 
        \sample_4[8]\, sample_4(7) => \sample_4[7]\, sample_4(6)
         => \sample_4[6]\, sample_4(5) => \sample_4[5]\, 
        sample_4(4) => \sample_4[4]\, sample_4(3) => 
        \sample_4[3]\, sample_4(2) => \sample_4[2]\, sample_4(1)
         => \sample_4[1]\, sample_4(0) => \sample_4[0]\, 
        sample_5(15) => \sample_5[15]\, sample_5(14) => 
        \sample_5[14]\, sample_5(13) => \sample_5[13]\, 
        sample_5(12) => \sample_5[12]\, sample_5(11) => 
        \sample_5[11]\, sample_5(10) => \sample_5[10]\, 
        sample_5(9) => \sample_5[9]\, sample_5(8) => 
        \sample_5[8]\, sample_5(7) => \sample_5[7]\, sample_5(6)
         => \sample_5[6]\, sample_5(5) => \sample_5[5]\, 
        sample_5(4) => \sample_5[4]\, sample_5(3) => 
        \sample_5[3]\, sample_5(2) => \sample_5[2]\, sample_5(1)
         => \sample_5[1]\, sample_5(0) => \sample_5[0]\, sdo_c(7)
         => sdo_c(7), sdo_c(6) => sdo_c(6), sdo_c(5) => sdo_c(5), 
        sdo_c(4) => sdo_c(4), sdo_c(3) => sdo_c(3), sdo_c(2) => 
        sdo_c(2), sdo_c(1) => sdo_c(1), sdo_c(0) => sdo_c(0), 
        sample_6(15) => \sample_6[15]\, sample_6(14) => 
        \sample_6[14]\, sample_6(13) => \sample_6[13]\, 
        sample_6(12) => \sample_6[12]\, sample_6(11) => 
        \sample_6[11]\, sample_6(10) => \sample_6[10]\, 
        sample_6(9) => \sample_6[9]\, sample_6(8) => 
        \sample_6[8]\, sample_6(7) => \sample_6[7]\, sample_6(6)
         => \sample_6[6]\, sample_6(5) => \sample_6[5]\, 
        sample_6(4) => \sample_6[4]\, sample_6(3) => 
        \sample_6[3]\, sample_6(2) => \sample_6[2]\, sample_6(1)
         => \sample_6[1]\, sample_6(0) => \sample_6[0]\, 
        cnv_rstn_c => cnv_rstn_c, cnv_clk_c => cnv_clk_c, cnv_c
         => cnv_c, sample_val => sample_val, sck_c => sck_c, 
        cnv_run_c => cnv_run_c, HRESETn_c => HRESETn_c, HCLK_c
         => HCLK_c);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out_RNO[97]\ : 
        MX2
      port map(A => \sample_filter_v2_out[97]\, B => 
        \sample_data_shaping_f2_f1_s[10]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_257[97]\);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[96]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_281[96]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[96]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I20_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[139]\, B => 
        \sample_filter_v2_out[121]\, Y => N187);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I19_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[122]\, B => 
        \sample_filter_v2_out[140]\, Y => N186);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[62]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[62]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[62]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I43_Y : 
        XA1A
      port map(A => \sample_filter_v2_out[104]\, B => 
        \sample_filter_v2_out[122]\, C => N187_0, Y => N275_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I48_Y : 
        NOR2
      port map(A => N255, B => N212_0, Y => N229_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I35_Y : 
        XAI1A
      port map(A => \sample_filter_v2_out[113]\, B => 
        \sample_filter_v2_out[131]\, C => N201, Y => N255);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I41_Y : 
        NOR2B
      port map(A => N191, B => N189, Y => N220_0);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[42]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[42]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[42]\);
    
    \SampleLoop_data_shaping.0.sample_data_shaping_out[71]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[71]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[71]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I27_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[132]\, B => 
        \sample_filter_v2_out[114]\, Y => N201);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I17_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[106]\, B => 
        \sample_filter_v2_out[124]\, Y => N182);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[52]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[52]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[52]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I30_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[111]\, B => 
        \sample_filter_v2_out[93]\, Y => N207);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[34]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[34]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[34]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I56_un1_Y : 
        OR3C
      port map(A => N275_0, B => N220, C => N278_0, Y => 
        I56_un1_Y);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I64_un1_Y : 
        OR2B
      port map(A => N268_0, B => N245, Y => I64_un1_Y);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I25_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[98]\, B => 
        \sample_filter_v2_out[116]\, Y => N198);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I25_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[116]\, B => 
        \sample_filter_v2_out[134]\, Y => N198_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I27_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[114]\, B => 
        \sample_filter_v2_out[132]\, Y => N202);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[111]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_349[111]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[111]\);
    
    \SampleLoop_data_shaping.8.sample_data_shaping_out[9]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[9]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[9]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I105_Y_0 : 
        AX1D
      port map(A => SUB_16x16_medium_area_I87_un1_Y, B => N202_0, 
        C => N203, Y => \sample_data_shaping_f2_f1_s[12]\);
    
    \SampleLoop_data_shaping.10.sample_data_shaping_out[7]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[7]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[7]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[48]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[48]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[48]\);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out[132]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[132]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[132]\);
    
    \SampleLoop_data_shaping.4.sample_data_shaping_out[31]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[31]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[31]\);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[16]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[16]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[16]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I33_Y : 
        NOR2B
      port map(A => N207, B => N205_0, Y => N212);
    
    \SampleLoop_data_shaping.11.sample_data_shaping_out_RNO[114]\ : 
        MX2
      port map(A => \sample_filter_v2_out[114]\, B => 
        \sample_data_shaping_f1_f0_s[11]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_277[114]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I86_un1_Y : 
        OA1
      port map(A => I71_un1_Y, B => N254, C => N205_0, Y => 
        I86_un1_Y);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out_RNO[113]\ : 
        MX2
      port map(A => \sample_filter_v2_out[113]\, B => 
        \sample_data_shaping_f1_f0_s[12]\, S => data_shaping_SP0, 
        Y => \sample_data_shaping_out_301[113]\);
    
    \SampleLoop_data_shaping.3.sample_data_shaping_out[50]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[50]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[50]\);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out_RNO[94]\ : 
        MX2
      port map(A => \sample_filter_v2_out[94]\, B => 
        \sample_data_shaping_f2_f1_s[13]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_329[94]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[2]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[2]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[2]\);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[66]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[66]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[66]\);
    
    \SampleLoop_data_shaping.1.sample_data_shaping_out[124]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_37[124]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[124]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I19_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[104]\, B => 
        \sample_filter_v2_out[122]\, Y => N186_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I25_S_0 : 
        XNOR2
      port map(A => \sample_filter_v2_out[134]\, B => 
        \sample_filter_v2_out[116]\, Y => N197);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I56_Y : 
        OR2B
      port map(A => SUB_16x16_medium_area_I56_Y_1, B => I56_un1_Y, 
        Y => N268_0);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[5]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[5]\, CLK => HCLK_c, CLR
         => HRESETn_c, Q => \sample_data_shaping_out[5]\);
    
    \SampleLoop_data_shaping.2.sample_data_shaping_out[105]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_65[105]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[105]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I104_Y_0 : 
        AX1A
      port map(A => N244, B => I64_un1_Y, C => N201_0, Y => 
        \sample_data_shaping_f2_f1_s[11]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[92]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_377[92]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[92]\);
    
    
        sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I89_un1_Y : 
        NOR2B
      port map(A => N268_0, B => N193, Y => 
        SUB_16x16_medium_area_I89_un1_Y);
    
    \SampleLoop_data_shaping.9.sample_data_shaping_out[44]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[44]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[44]\);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I56_Y_0 : 
        AO18
      port map(A => N190_0, B => \sample_filter_v2_out[137]\, C
         => \sample_filter_v2_out[119]\, Y => 
        SUB_16x16_medium_area_I56_Y_0_0);
    
    \SampleLoop_data_shaping.14.sample_data_shaping_out[21]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[21]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[21]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I35_Y : 
        NOR2B
      port map(A => N203, B => N201_0, Y => N255_0);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out[38]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[38]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[38]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I56_Y_1 : 
        AOI1B
      port map(A => N274, B => N220, C => 
        SUB_16x16_medium_area_I56_Y_0, Y => 
        SUB_16x16_medium_area_I56_Y_1);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I50_Y : 
        NOR2B
      port map(A => N265_0, B => N216_0, Y => N245);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I56_un1_Y_0 : 
        NOR2B
      port map(A => N220_0, B => N275, Y => 
        SUB_16x16_medium_area_I56_un1_Y_0);
    
    \SampleLoop_data_shaping.7.sample_data_shaping_out[100]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_185[100]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[100]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I98_Y_0 : 
        XOR2
      port map(A => N280, B => N189_0, Y => 
        \sample_data_shaping_f2_f1_s[5]\);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[95]\ : 
        DFN1C0
      port map(D => \sample_data_shaping_out_305[95]\, CLK => 
        HCLK_c, CLR => HRESETn_c, Q => 
        \sample_data_shaping_out[95]\);
    
    \SampleLoop_data_shaping.6.sample_data_shaping_out[65]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[65]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[65]\);
    
    \SampleLoop_data_shaping.15.sample_data_shaping_out_RNO[92]\ : 
        MX2
      port map(A => \sample_filter_v2_out[92]\, B => 
        \sample_data_shaping_f2_f1_s[15]\, S => data_shaping_SP1, 
        Y => \sample_data_shaping_out_377[92]\);
    
    \SampleLoop_data_shaping.12.sample_data_shaping_out[131]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[131]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[131]\);
    
    \SampleLoop_data_shaping.13.sample_data_shaping_out[22]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[22]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[22]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I91_un1_Y : 
        NOR2B
      port map(A => N278, B => N185, Y => 
        SUB_16x16_medium_area_I91_un1_Y);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I53_Y_0 : 
        AO18
      port map(A => N182_0, B => \sample_filter_v2_out[141]\, C
         => \sample_filter_v2_out[123]\, Y => 
        SUB_16x16_medium_area_I53_Y_0_0);
    
    \SampleLoop_data_shaping.5.sample_data_shaping_out[12]\ : 
        DFN1C0
      port map(D => \sample_filter_v2_out[12]\, CLK => HCLK_c, 
        CLR => HRESETn_c, Q => \sample_data_shaping_out[12]\);
    
    sample_data_shaping_f2_f1_s_0_0_SUB_16x16_medium_area_I23_CO1 : 
        NOR2A
      port map(A => \sample_filter_v2_out[100]\, B => 
        \sample_filter_v2_out[118]\, Y => N194_0);
    
    sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I97_Y_0 : 
        AX1D
      port map(A => SUB_16x16_medium_area_I91_un1_Y, B => N186, C
         => N187, Y => \sample_data_shaping_f1_f0_s[4]\);
    
    
        sample_data_shaping_f1_f0_s_0_0_SUB_16x16_medium_area_I100_Y_0 : 
        XNOR3
      port map(A => \sample_filter_v2_out[118]\, B => 
        \sample_filter_v2_out[136]\, C => N268, Y => 
        \sample_data_shaping_f1_f0_s[7]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity lpp_top_lfr_wf_picker is

    port( cnv_run         : in    std_logic;
          cnv             : out   std_logic;
          sck             : out   std_logic;
          sdo             : in    std_logic_vector(7 downto 0);
          cnv_clk         : in    std_logic;
          cnv_rstn        : in    std_logic;
          HCLK            : in    std_logic;
          HRESETn         : in    std_logic;
          apbi            : in    std_logic_vector(121 downto 0);
          apbo            : out   std_logic_vector(131 downto 0);
          AHB_Master_In   : in    std_logic_vector(90 downto 0);
          AHB_Master_Out  : out   std_logic_vector(370 downto 0);
          coarse_time_0   : in    std_logic;
          data_shaping_BW : out   std_logic
        );

end lpp_top_lfr_wf_picker;

architecture DEF_ARCH of lpp_top_lfr_wf_picker is 

  component OUTBUF
    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component INBUF
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component lpp_top_apbreg
    port( status_full_ack    : out   std_logic_vector(3 downto 0);
          prdata_c           : out   std_logic_vector(31 downto 0);
          pirq_c             : out   std_logic_vector(15 to 15);
          addr_data_f2       : out   std_logic_vector(31 downto 0);
          status_new_err_3   : in    std_logic := 'U';
          status_new_err_0_2 : in    std_logic := 'U';
          status_new_err_0_0 : in    std_logic := 'U';
          status_new_err_0_1 : in    std_logic := 'U';
          status_full_err_0  : in    std_logic_vector(3 downto 0) := (others => 'U');
          status_full        : in    std_logic_vector(3 downto 0) := (others => 'U');
          addr_data_f3       : out   std_logic_vector(31 downto 0);
          nb_burst_available : out   std_logic_vector(10 downto 0);
          addr_data_f1       : out   std_logic_vector(31 downto 0);
          delta_f2_f1        : out   std_logic_vector(9 downto 0);
          addr_data_f0       : out   std_logic_vector(31 downto 0);
          delta_f2_f0        : out   std_logic_vector(9 downto 0);
          delta_snapshot     : out   std_logic_vector(15 downto 0);
          nb_snapshot_param  : out   std_logic_vector(10 downto 0);
          apbi_c_81          : in    std_logic := 'U';
          apbi_c_80          : in    std_logic := 'U';
          apbi_c_79          : in    std_logic := 'U';
          apbi_c_78          : in    std_logic := 'U';
          apbi_c_77          : in    std_logic := 'U';
          apbi_c_76          : in    std_logic := 'U';
          apbi_c_75          : in    std_logic := 'U';
          apbi_c_74          : in    std_logic := 'U';
          apbi_c_73          : in    std_logic := 'U';
          apbi_c_72          : in    std_logic := 'U';
          apbi_c_71          : in    std_logic := 'U';
          apbi_c_70          : in    std_logic := 'U';
          apbi_c_69          : in    std_logic := 'U';
          apbi_c_68          : in    std_logic := 'U';
          apbi_c_67          : in    std_logic := 'U';
          apbi_c_66          : in    std_logic := 'U';
          apbi_c_65          : in    std_logic := 'U';
          apbi_c_64          : in    std_logic := 'U';
          apbi_c_63          : in    std_logic := 'U';
          apbi_c_62          : in    std_logic := 'U';
          apbi_c_61          : in    std_logic := 'U';
          apbi_c_60          : in    std_logic := 'U';
          apbi_c_59          : in    std_logic := 'U';
          apbi_c_58          : in    std_logic := 'U';
          apbi_c_57          : in    std_logic := 'U';
          apbi_c_56          : in    std_logic := 'U';
          apbi_c_55          : in    std_logic := 'U';
          apbi_c_24          : in    std_logic := 'U';
          apbi_c_23          : in    std_logic := 'U';
          apbi_c_0           : in    std_logic := 'U';
          apbi_c_50          : in    std_logic := 'U';
          apbi_c_51          : in    std_logic := 'U';
          apbi_c_52          : in    std_logic := 'U';
          apbi_c_16          : in    std_logic := 'U';
          apbi_c_49          : in    std_logic := 'U';
          apbi_c_22          : in    std_logic := 'U';
          apbi_c_20          : in    std_logic := 'U';
          apbi_c_19          : in    std_logic := 'U';
          apbi_c_21          : in    std_logic := 'U';
          apbi_c_54          : in    std_logic := 'U';
          apbi_c_53          : in    std_logic := 'U';
          data_shaping_R0    : out   std_logic;
          data_shaping_R1    : out   std_logic;
          enable_f0          : out   std_logic;
          data_shaping_BW_c  : out   std_logic;
          burst_f2           : out   std_logic;
          burst_f1           : out   std_logic;
          burst_f0           : out   std_logic;
          enable_f3          : out   std_logic;
          enable_f2          : out   std_logic;
          data_shaping_SP1   : out   std_logic;
          enable_f1          : out   std_logic;
          data_shaping_SP0   : out   std_logic;
          data_shaping_R1_0  : out   std_logic;
          HRESETn_c          : in    std_logic := 'U';
          HCLK_c             : in    std_logic := 'U';
          data_shaping_R0_0  : out   std_logic
        );
  end component;

  component lpp_top_lfr_wf_picker_ip
    port( nb_snapshot_param            : in    std_logic_vector(10 downto 0) := (others => 'U');
          delta_f2_f0                  : in    std_logic_vector(9 downto 0) := (others => 'U');
          delta_snapshot               : in    std_logic_vector(15 downto 0) := (others => 'U');
          delta_f2_f1                  : in    std_logic_vector(9 downto 0) := (others => 'U');
          status_new_err               : out   std_logic_vector(3 downto 0);
          hwdata_c                     : out   std_logic_vector(31 downto 0);
          addr_data_f0                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f1                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f2                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          addr_data_f3                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          status_full                  : out   std_logic_vector(3 downto 0);
          status_full_err              : out   std_logic_vector(3 downto 0);
          nb_burst_available           : in    std_logic_vector(10 downto 0) := (others => 'U');
          haddr_c                      : out   std_logic_vector(31 downto 0);
          AHB_Master_In_c_3            : in    std_logic := 'U';
          AHB_Master_In_c_0            : in    std_logic := 'U';
          AHB_Master_In_c_4            : in    std_logic := 'U';
          AHB_Master_In_c_5            : in    std_logic := 'U';
          hsize_c                      : out   std_logic_vector(1 downto 0);
          htrans_c                     : out   std_logic_vector(1 downto 0);
          hburst_c                     : out   std_logic_vector(2 downto 0);
          status_full_ack              : in    std_logic_vector(3 downto 0) := (others => 'U');
          sdo_c                        : in    std_logic_vector(7 downto 0) := (others => 'U');
          coarse_time_0_c              : in    std_logic := 'U';
          enable_f0                    : in    std_logic := 'U';
          data_shaping_R0              : in    std_logic := 'U';
          data_shaping_R0_0            : in    std_logic := 'U';
          burst_f0                     : in    std_logic := 'U';
          data_shaping_R1              : in    std_logic := 'U';
          data_shaping_R1_0            : in    std_logic := 'U';
          enable_f1                    : in    std_logic := 'U';
          burst_f1                     : in    std_logic := 'U';
          enable_f2                    : in    std_logic := 'U';
          burst_f2                     : in    std_logic := 'U';
          enable_f3                    : in    std_logic := 'U';
          N_43                         : out   std_logic;
          IdlePhase_RNI03G71           : out   std_logic;
          hwrite_c                     : out   std_logic;
          lpp_top_lfr_wf_picker_ip_GND : in    std_logic := 'U';
          lpp_top_lfr_wf_picker_ip_VCC : in    std_logic := 'U';
          cnv_run_c                    : in    std_logic := 'U';
          sck_c                        : out   std_logic;
          cnv_c                        : out   std_logic;
          cnv_clk_c                    : in    std_logic := 'U';
          cnv_rstn_c                   : in    std_logic := 'U';
          data_shaping_SP0             : in    std_logic := 'U';
          data_shaping_SP1             : in    std_logic := 'U';
          HRESETn_c                    : in    std_logic := 'U';
          HCLK_c                       : in    std_logic := 'U'
        );
  end component;

  component CLKBUF
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

    signal \status_full[0]\, \status_full[1]\, \status_full[2]\, 
        \status_full[3]\, \status_full_ack[0]\, 
        \status_full_ack[1]\, \status_full_ack[2]\, 
        \status_full_ack[3]\, \status_full_err[0]\, 
        \status_full_err[1]\, \status_full_err[2]\, 
        \status_full_err[3]\, \status_new_err[0]\, 
        \status_new_err[1]\, \status_new_err[2]\, 
        \status_new_err[3]\, data_shaping_SP0, data_shaping_SP1, 
        data_shaping_R0, data_shaping_R1, \delta_snapshot[0]\, 
        \delta_snapshot[1]\, \delta_snapshot[2]\, 
        \delta_snapshot[3]\, \delta_snapshot[4]\, 
        \delta_snapshot[5]\, \delta_snapshot[6]\, 
        \delta_snapshot[7]\, \delta_snapshot[8]\, 
        \delta_snapshot[9]\, \delta_snapshot[10]\, 
        \delta_snapshot[11]\, \delta_snapshot[12]\, 
        \delta_snapshot[13]\, \delta_snapshot[14]\, 
        \delta_snapshot[15]\, \delta_f2_f1[0]\, \delta_f2_f1[1]\, 
        \delta_f2_f1[2]\, \delta_f2_f1[3]\, \delta_f2_f1[4]\, 
        \delta_f2_f1[5]\, \delta_f2_f1[6]\, \delta_f2_f1[7]\, 
        \delta_f2_f1[8]\, \delta_f2_f1[9]\, \delta_f2_f0[0]\, 
        \delta_f2_f0[1]\, \delta_f2_f0[2]\, \delta_f2_f0[3]\, 
        \delta_f2_f0[4]\, \delta_f2_f0[5]\, \delta_f2_f0[6]\, 
        \delta_f2_f0[7]\, \delta_f2_f0[8]\, \delta_f2_f0[9]\, 
        \nb_burst_available[0]\, \nb_burst_available[1]\, 
        \nb_burst_available[2]\, \nb_burst_available[3]\, 
        \nb_burst_available[4]\, \nb_burst_available[5]\, 
        \nb_burst_available[6]\, \nb_burst_available[7]\, 
        \nb_burst_available[8]\, \nb_burst_available[9]\, 
        \nb_burst_available[10]\, \nb_snapshot_param[0]\, 
        \nb_snapshot_param[1]\, \nb_snapshot_param[2]\, 
        \nb_snapshot_param[3]\, \nb_snapshot_param[4]\, 
        \nb_snapshot_param[5]\, \nb_snapshot_param[6]\, 
        \nb_snapshot_param[7]\, \nb_snapshot_param[8]\, 
        \nb_snapshot_param[9]\, \nb_snapshot_param[10]\, 
        enable_f0, enable_f1, enable_f2, enable_f3, burst_f0, 
        burst_f1, burst_f2, \addr_data_f0[0]\, \addr_data_f0[1]\, 
        \addr_data_f0[2]\, \addr_data_f0[3]\, \addr_data_f0[4]\, 
        \addr_data_f0[5]\, \addr_data_f0[6]\, \addr_data_f0[7]\, 
        \addr_data_f0[8]\, \addr_data_f0[9]\, \addr_data_f0[10]\, 
        \addr_data_f0[11]\, \addr_data_f0[12]\, 
        \addr_data_f0[13]\, \addr_data_f0[14]\, 
        \addr_data_f0[15]\, \addr_data_f0[16]\, 
        \addr_data_f0[17]\, \addr_data_f0[18]\, 
        \addr_data_f0[19]\, \addr_data_f0[20]\, 
        \addr_data_f0[21]\, \addr_data_f0[22]\, 
        \addr_data_f0[23]\, \addr_data_f0[24]\, 
        \addr_data_f0[25]\, \addr_data_f0[26]\, 
        \addr_data_f0[27]\, \addr_data_f0[28]\, 
        \addr_data_f0[29]\, \addr_data_f0[30]\, 
        \addr_data_f0[31]\, \addr_data_f1[0]\, \addr_data_f1[1]\, 
        \addr_data_f1[2]\, \addr_data_f1[3]\, \addr_data_f1[4]\, 
        \addr_data_f1[5]\, \addr_data_f1[6]\, \addr_data_f1[7]\, 
        \addr_data_f1[8]\, \addr_data_f1[9]\, \addr_data_f1[10]\, 
        \addr_data_f1[11]\, \addr_data_f1[12]\, 
        \addr_data_f1[13]\, \addr_data_f1[14]\, 
        \addr_data_f1[15]\, \addr_data_f1[16]\, 
        \addr_data_f1[17]\, \addr_data_f1[18]\, 
        \addr_data_f1[19]\, \addr_data_f1[20]\, 
        \addr_data_f1[21]\, \addr_data_f1[22]\, 
        \addr_data_f1[23]\, \addr_data_f1[24]\, 
        \addr_data_f1[25]\, \addr_data_f1[26]\, 
        \addr_data_f1[27]\, \addr_data_f1[28]\, 
        \addr_data_f1[29]\, \addr_data_f1[30]\, 
        \addr_data_f1[31]\, \addr_data_f2[0]\, \addr_data_f2[1]\, 
        \addr_data_f2[2]\, \addr_data_f2[3]\, \addr_data_f2[4]\, 
        \addr_data_f2[5]\, \addr_data_f2[6]\, \addr_data_f2[7]\, 
        \addr_data_f2[8]\, \addr_data_f2[9]\, \addr_data_f2[10]\, 
        \addr_data_f2[11]\, \addr_data_f2[12]\, 
        \addr_data_f2[13]\, \addr_data_f2[14]\, 
        \addr_data_f2[15]\, \addr_data_f2[16]\, 
        \addr_data_f2[17]\, \addr_data_f2[18]\, 
        \addr_data_f2[19]\, \addr_data_f2[20]\, 
        \addr_data_f2[21]\, \addr_data_f2[22]\, 
        \addr_data_f2[23]\, \addr_data_f2[24]\, 
        \addr_data_f2[25]\, \addr_data_f2[26]\, 
        \addr_data_f2[27]\, \addr_data_f2[28]\, 
        \addr_data_f2[29]\, \addr_data_f2[30]\, 
        \addr_data_f2[31]\, \addr_data_f3[0]\, \addr_data_f3[1]\, 
        \addr_data_f3[2]\, \addr_data_f3[3]\, \addr_data_f3[4]\, 
        \addr_data_f3[5]\, \addr_data_f3[6]\, \addr_data_f3[7]\, 
        \addr_data_f3[8]\, \addr_data_f3[9]\, \addr_data_f3[10]\, 
        \addr_data_f3[11]\, \addr_data_f3[12]\, 
        \addr_data_f3[13]\, \addr_data_f3[14]\, 
        \addr_data_f3[15]\, \addr_data_f3[16]\, 
        \addr_data_f3[17]\, \addr_data_f3[18]\, 
        \addr_data_f3[19]\, \addr_data_f3[20]\, 
        \addr_data_f3[21]\, \addr_data_f3[22]\, 
        \addr_data_f3[23]\, \addr_data_f3[24]\, 
        \addr_data_f3[25]\, \addr_data_f3[26]\, 
        \addr_data_f3[27]\, \addr_data_f3[28]\, 
        \addr_data_f3[29]\, \addr_data_f3[30]\, 
        \addr_data_f3[31]\, IdlePhase_RNI03G71, 
        \lpp_top_lfr_wf_picker_ip_1.lpp_waveform_1.pp_waveform_dma_1.DMA2AHB_1.N_43\, 
        cnv_run_c, cnv_c, sck_c, \sdo_c[0]\, \sdo_c[1]\, 
        \sdo_c[2]\, \sdo_c[3]\, \sdo_c[4]\, \sdo_c[5]\, 
        \sdo_c[6]\, \sdo_c[7]\, cnv_clk_c, cnv_rstn_c, HCLK_c, 
        HRESETn_c, \apbi_c[0]\, \apbi_c[16]\, \apbi_c[19]\, 
        \apbi_c[20]\, \apbi_c[21]\, \apbi_c[22]\, \apbi_c[23]\, 
        \apbi_c[24]\, \apbi_c[49]\, \apbi_c[50]\, \apbi_c[51]\, 
        \apbi_c[52]\, \apbi_c[53]\, \apbi_c[54]\, \apbi_c[55]\, 
        \apbi_c[56]\, \apbi_c[57]\, \apbi_c[58]\, \apbi_c[59]\, 
        \apbi_c[60]\, \apbi_c[61]\, \apbi_c[62]\, \apbi_c[63]\, 
        \apbi_c[64]\, \apbi_c[65]\, \apbi_c[66]\, \apbi_c[67]\, 
        \apbi_c[68]\, \apbi_c[69]\, \apbi_c[70]\, \apbi_c[71]\, 
        \apbi_c[72]\, \apbi_c[73]\, \apbi_c[74]\, \apbi_c[75]\, 
        \apbi_c[76]\, \apbi_c[77]\, \apbi_c[78]\, \apbi_c[79]\, 
        \apbi_c[80]\, \apbi_c[81]\, \apbo.prdata_c[0]\, 
        \apbo.prdata_c[1]\, \apbo.prdata_c[2]\, 
        \apbo.prdata_c[3]\, \apbo.prdata_c[4]\, 
        \apbo.prdata_c[5]\, \apbo.prdata_c[6]\, 
        \apbo.prdata_c[7]\, \apbo.prdata_c[8]\, 
        \apbo.prdata_c[9]\, \apbo.prdata_c[10]\, 
        \apbo.prdata_c[11]\, \apbo.prdata_c[12]\, 
        \apbo.prdata_c[13]\, \apbo.prdata_c[14]\, 
        \apbo.prdata_c[15]\, \apbo.prdata_c[16]\, 
        \apbo.prdata_c[17]\, \apbo.prdata_c[18]\, 
        \apbo.prdata_c[19]\, \apbo.prdata_c[20]\, 
        \apbo.prdata_c[21]\, \apbo.prdata_c[22]\, 
        \apbo.prdata_c[23]\, \apbo.prdata_c[24]\, 
        \apbo.prdata_c[25]\, \apbo.prdata_c[26]\, 
        \apbo.prdata_c[27]\, \apbo.prdata_c[28]\, 
        \apbo.prdata_c[29]\, \apbo.prdata_c[30]\, 
        \apbo.prdata_c[31]\, \apbo.pirq_c[15]\, 
        \AHB_Master_In_c[13]\, \AHB_Master_In_c[16]\, 
        \AHB_Master_In_c[17]\, \AHB_Master_In_c[18]\, 
        \AHB_Master_Out.htrans_c[0]\, 
        \AHB_Master_Out.htrans_c[1]\, \AHB_Master_Out.haddr_c[0]\, 
        \AHB_Master_Out.haddr_c[1]\, \AHB_Master_Out.haddr_c[2]\, 
        \AHB_Master_Out.haddr_c[3]\, \AHB_Master_Out.haddr_c[4]\, 
        \AHB_Master_Out.haddr_c[5]\, \AHB_Master_Out.haddr_c[6]\, 
        \AHB_Master_Out.haddr_c[7]\, \AHB_Master_Out.haddr_c[8]\, 
        \AHB_Master_Out.haddr_c[9]\, \AHB_Master_Out.haddr_c[10]\, 
        \AHB_Master_Out.haddr_c[11]\, 
        \AHB_Master_Out.haddr_c[12]\, 
        \AHB_Master_Out.haddr_c[13]\, 
        \AHB_Master_Out.haddr_c[14]\, 
        \AHB_Master_Out.haddr_c[15]\, 
        \AHB_Master_Out.haddr_c[16]\, 
        \AHB_Master_Out.haddr_c[17]\, 
        \AHB_Master_Out.haddr_c[18]\, 
        \AHB_Master_Out.haddr_c[19]\, 
        \AHB_Master_Out.haddr_c[20]\, 
        \AHB_Master_Out.haddr_c[21]\, 
        \AHB_Master_Out.haddr_c[22]\, 
        \AHB_Master_Out.haddr_c[23]\, 
        \AHB_Master_Out.haddr_c[24]\, 
        \AHB_Master_Out.haddr_c[25]\, 
        \AHB_Master_Out.haddr_c[26]\, 
        \AHB_Master_Out.haddr_c[27]\, 
        \AHB_Master_Out.haddr_c[28]\, 
        \AHB_Master_Out.haddr_c[29]\, 
        \AHB_Master_Out.haddr_c[30]\, 
        \AHB_Master_Out.haddr_c[31]\, \AHB_Master_Out.hwrite_c\, 
        \AHB_Master_Out.hsize_c[0]\, \AHB_Master_Out.hsize_c[1]\, 
        \AHB_Master_Out.hburst_c[0]\, 
        \AHB_Master_Out.hburst_c[1]\, 
        \AHB_Master_Out.hburst_c[2]\, 
        \AHB_Master_Out.hwdata_c[0]\, 
        \AHB_Master_Out.hwdata_c[1]\, 
        \AHB_Master_Out.hwdata_c[2]\, 
        \AHB_Master_Out.hwdata_c[3]\, 
        \AHB_Master_Out.hwdata_c[4]\, 
        \AHB_Master_Out.hwdata_c[5]\, 
        \AHB_Master_Out.hwdata_c[6]\, 
        \AHB_Master_Out.hwdata_c[7]\, 
        \AHB_Master_Out.hwdata_c[8]\, 
        \AHB_Master_Out.hwdata_c[9]\, 
        \AHB_Master_Out.hwdata_c[10]\, 
        \AHB_Master_Out.hwdata_c[11]\, 
        \AHB_Master_Out.hwdata_c[12]\, 
        \AHB_Master_Out.hwdata_c[13]\, 
        \AHB_Master_Out.hwdata_c[14]\, 
        \AHB_Master_Out.hwdata_c[15]\, 
        \AHB_Master_Out.hwdata_c[16]\, 
        \AHB_Master_Out.hwdata_c[17]\, 
        \AHB_Master_Out.hwdata_c[18]\, 
        \AHB_Master_Out.hwdata_c[19]\, 
        \AHB_Master_Out.hwdata_c[20]\, 
        \AHB_Master_Out.hwdata_c[21]\, 
        \AHB_Master_Out.hwdata_c[22]\, 
        \AHB_Master_Out.hwdata_c[23]\, 
        \AHB_Master_Out.hwdata_c[24]\, 
        \AHB_Master_Out.hwdata_c[25]\, 
        \AHB_Master_Out.hwdata_c[26]\, 
        \AHB_Master_Out.hwdata_c[27]\, 
        \AHB_Master_Out.hwdata_c[28]\, 
        \AHB_Master_Out.hwdata_c[29]\, 
        \AHB_Master_Out.hwdata_c[30]\, 
        \AHB_Master_Out.hwdata_c[31]\, \VCC\, \GND\, 
        coarse_time_0_c, data_shaping_BW_c, data_shaping_R1_0, 
        data_shaping_R0_0, GND_0, VCC_0 : std_logic;

    for all : lpp_top_apbreg
	Use entity work.lpp_top_apbreg(DEF_ARCH);
    for all : lpp_top_lfr_wf_picker_ip
	Use entity work.lpp_top_lfr_wf_picker_ip(DEF_ARCH);
begin 


    \apbo_pad[90]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(90));
    
    \apbi_pad[78]\ : INBUF
      port map(PAD => apbi(78), Y => \apbi_c[78]\);
    
    \apbo_pad[113]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(113));
    
    \AHB_Master_Out_pad[189]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(189));
    
    \AHB_Master_Out_pad[170]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(170));
    
    \apbo_pad[106]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(106));
    
    \apbi_pad[23]\ : INBUF
      port map(PAD => apbi(23), Y => \apbi_c[23]\);
    
    \apbo_pad[18]\ : OUTBUF
      port map(D => \apbo.prdata_c[18]\, PAD => apbo(18));
    
    \AHB_Master_Out_pad[15]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[11]\, PAD => 
        AHB_Master_Out(15));
    
    \AHB_Master_Out_pad[6]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[2]\, PAD => 
        AHB_Master_Out(6));
    
    \AHB_Master_Out_pad[4]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[0]\, PAD => 
        AHB_Master_Out(4));
    
    \AHB_Master_Out_pad[40]\ : OUTBUF
      port map(D => \AHB_Master_Out.hburst_c[0]\, PAD => 
        AHB_Master_Out(40));
    
    \AHB_Master_Out_pad[176]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(176));
    
    \AHB_Master_Out_pad[132]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(132));
    
    \AHB_Master_Out_pad[51]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[4]\, PAD => 
        AHB_Master_Out(51));
    
    \apbo_pad[102]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(102));
    
    \AHB_Master_Out_pad[257]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(257));
    
    \apbo_pad[124]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(124));
    
    \AHB_Master_Out_pad[318]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(318));
    
    \apbo_pad[91]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(91));
    
    \AHB_Master_Out_pad[328]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(328));
    
    \AHB_Master_In_pad[17]\ : INBUF
      port map(PAD => AHB_Master_In(17), Y => 
        \AHB_Master_In_c[17]\);
    
    \apbo_pad[95]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(95));
    
    \AHB_Master_Out_pad[348]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(348));
    
    \AHB_Master_Out_pad[259]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(259));
    
    \AHB_Master_Out_pad[332]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(332));
    
    \AHB_Master_Out_pad[12]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[8]\, PAD => 
        AHB_Master_Out(12));
    
    \AHB_Master_Out_pad[1]\ : OUTBUF
      port map(D => 
        \lpp_top_lfr_wf_picker_ip_1.lpp_waveform_1.pp_waveform_dma_1.DMA2AHB_1.N_43\, 
        PAD => AHB_Master_Out(1));
    
    \sdo_pad[4]\ : INBUF
      port map(PAD => sdo(4), Y => \sdo_c[4]\);
    
    \AHB_Master_Out_pad[46]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(46));
    
    \apbo_pad[48]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(48));
    
    \AHB_Master_Out_pad[214]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(214));
    
    \apbo_pad[6]\ : OUTBUF
      port map(D => \apbo.prdata_c[6]\, PAD => apbo(6));
    
    \AHB_Master_Out_pad[224]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(224));
    
    \AHB_Master_Out_pad[244]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(244));
    
    \AHB_Master_Out_pad[150]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(150));
    
    \AHB_Master_Out_pad[368]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(368));
    
    \AHB_Master_Out_pad[339]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(339));
    
    \AHB_Master_Out_pad[297]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(297));
    
    \AHB_Master_Out_pad[201]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(201));
    
    \AHB_Master_Out_pad[47]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[0]\, PAD => 
        AHB_Master_Out(47));
    
    \AHB_Master_Out_pad[307]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(307));
    
    \AHB_Master_Out_pad[213]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(213));
    
    \apbo_pad[57]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(57));
    
    \AHB_Master_Out_pad[223]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(223));
    
    \AHB_Master_Out_pad[156]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(156));
    
    \AHB_Master_Out_pad[111]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(111));
    
    \apbi_pad[76]\ : INBUF
      port map(PAD => apbi(76), Y => \apbi_c[76]\);
    
    \AHB_Master_Out_pad[243]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(243));
    
    \AHB_Master_Out_pad[121]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(121));
    
    \apbo_pad[89]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(89));
    
    \AHB_Master_Out_pad[299]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(299));
    
    \AHB_Master_Out_pad[141]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(141));
    
    \AHB_Master_Out_pad[49]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[2]\, PAD => 
        AHB_Master_Out(49));
    
    \AHB_Master_Out_pad[182]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(182));
    
    \apbo_pad[16]\ : OUTBUF
      port map(D => \apbo.prdata_c[16]\, PAD => apbo(16));
    
    \AHB_Master_Out_pad[264]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(264));
    
    \AHB_Master_Out_pad[301]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(301));
    
    \apbo_pad[53]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(53));
    
    \AHB_Master_Out_pad[190]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(190));
    
    \AHB_Master_Out_pad[232]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(232));
    
    \AHB_Master_In_pad[16]\ : INBUF
      port map(PAD => AHB_Master_In(16), Y => 
        \AHB_Master_In_c[16]\);
    
    \AHB_Master_Out_pad[263]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(263));
    
    \AHB_Master_Out_pad[25]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[21]\, PAD => 
        AHB_Master_Out(25));
    
    \AHB_Master_Out_pad[161]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(161));
    
    \AHB_Master_Out_pad[196]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(196));
    
    \AHB_Master_Out_pad[134]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(134));
    
    \AHB_Master_Out_pad[0]\ : OUTBUF
      port map(D => IdlePhase_RNI03G71, PAD => AHB_Master_Out(0));
    
    \AHB_Master_In_pad[13]\ : INBUF
      port map(PAD => AHB_Master_In(13), Y => 
        \AHB_Master_In_c[13]\);
    
    sck_pad : OUTBUF
      port map(D => sck_c, PAD => sck);
    
    \apbi_pad[68]\ : INBUF
      port map(PAD => apbi(68), Y => \apbi_c[68]\);
    
    \AHB_Master_Out_pad[200]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(200));
    
    \AHB_Master_Out_pad[61]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[14]\, PAD => 
        AHB_Master_Out(61));
    
    \AHB_Master_Out_pad[105]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(105));
    
    \AHB_Master_Out_pad[117]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(117));
    
    \AHB_Master_Out_pad[127]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(127));
    
    \AHB_Master_Out_pad[147]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(147));
    
    \apbo_pad[46]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(46));
    
    \AHB_Master_Out_pad[335]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(335));
    
    \apbi_pad[74]\ : INBUF
      port map(PAD => apbi(74), Y => \apbi_c[74]\);
    
    \AHB_Master_Out_pad[22]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[18]\, PAD => 
        AHB_Master_Out(22));
    
    \apbo_pad[131]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(131));
    
    \apbo_pad[7]\ : OUTBUF
      port map(D => \apbo.prdata_c[7]\, PAD => apbo(7));
    
    \AHB_Master_Out_pad[206]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(206));
    
    coarse_time_0_pad : INBUF
      port map(PAD => coarse_time_0, Y => coarse_time_0_c);
    
    \apbo_pad[127]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(127));
    
    \apbo_pad[14]\ : OUTBUF
      port map(D => \apbo.prdata_c[14]\, PAD => apbo(14));
    
    \AHB_Master_Out_pad[108]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(108));
    
    \apbo_pad[119]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(119));
    
    \AHB_Master_Out_pad[167]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(167));
    
    \AHB_Master_Out_pad[14]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[10]\, PAD => 
        AHB_Master_Out(14));
    
    \AHB_Master_Out_pad[31]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[27]\, PAD => 
        AHB_Master_Out(31));
    
    \AHB_Master_Out_pad[282]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(282));
    
    \AHB_Master_Out_pad[184]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(184));
    
    \AHB_Master_Out_pad[133]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(133));
    
    \apbo_pad[98]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(98));
    
    \AHB_Master_Out_pad[303]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(303));
    
    \apbo_pad[44]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(44));
    
    \apbi_pad[66]\ : INBUF
      port map(PAD => apbi(66), Y => \apbi_c[66]\);
    
    \AHB_Master_Out_pad[274]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(274));
    
    \apbo_pad[79]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(79));
    
    \AHB_Master_Out_pad[211]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(211));
    
    \apbo_pad[32]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(32));
    
    \AHB_Master_Out_pad[317]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(317));
    
    \AHB_Master_Out_pad[221]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(221));
    
    \AHB_Master_Out_pad[327]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(327));
    
    \AHB_Master_Out_pad[241]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(241));
    
    \apbi_pad[52]\ : INBUF
      port map(PAD => apbi(52), Y => \apbi_c[52]\);
    
    \AHB_Master_Out_pad[347]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(347));
    
    \apbo_pad[22]\ : OUTBUF
      port map(D => \apbo.prdata_c[22]\, PAD => apbo(22));
    
    \AHB_Master_Out_pad[7]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[3]\, PAD => 
        AHB_Master_Out(7));
    
    \AHB_Master_Out_pad[336]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(336));
    
    \AHB_Master_Out_pad[273]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(273));
    
    \apbo_pad[116]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(116));
    
    \AHB_Master_Out_pad[171]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(171));
    
    \apbo_pad[108]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(108));
    
    \sdo_pad[1]\ : INBUF
      port map(PAD => sdo(1), Y => \sdo_c[1]\);
    
    \AHB_Master_Out_pad[98]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(98));
    
    \AHB_Master_Out_pad[13]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[9]\, PAD => 
        AHB_Master_Out(13));
    
    \AHB_Master_Out_pad[358]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(358));
    
    \AHB_Master_Out_pad[311]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(311));
    
    \apbo_pad[30]\ : OUTBUF
      port map(D => \apbo.prdata_c[30]\, PAD => apbo(30));
    
    \AHB_Master_Out_pad[321]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(321));
    
    \AHB_Master_Out_pad[208]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(208));
    
    \apbo_pad[62]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(62));
    
    \apbo_pad[112]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(112));
    
    \AHB_Master_Out_pad[341]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(341));
    
    \apbi_pad[50]\ : INBUF
      port map(PAD => apbi(50), Y => \apbi_c[50]\);
    
    \apbo_pad[20]\ : OUTBUF
      port map(D => \apbo.prdata_c[20]\, PAD => apbo(20));
    
    \AHB_Master_Out_pad[261]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(261));
    
    \AHB_Master_Out_pad[367]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(367));
    
    \AHB_Master_Out_pad[90]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(90));
    
    \AHB_Master_Out_pad[183]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(183));
    
    \AHB_Master_Out_pad[109]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(109));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \AHB_Master_Out_pad[45]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(45));
    
    \AHB_Master_Out_pad[254]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(254));
    
    \AHB_Master_Out_pad[210]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(210));
    
    \AHB_Master_Out_pad[220]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(220));
    
    \AHB_Master_Out_pad[115]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(115));
    
    \apbo_pad[60]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(60));
    
    \apbi_pad[77]\ : INBUF
      port map(PAD => apbi(77), Y => \apbi_c[77]\);
    
    \apbi_pad[64]\ : INBUF
      port map(PAD => apbi(64), Y => \apbi_c[64]\);
    
    \AHB_Master_Out_pad[240]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(240));
    
    \AHB_Master_Out_pad[125]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(125));
    
    \apbo_pad[96]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(96));
    
    \AHB_Master_Out_pad[145]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(145));
    
    \apbo_pad[31]\ : OUTBUF
      port map(D => \apbo.prdata_c[31]\, PAD => apbo(31));
    
    \AHB_Master_Out_pad[361]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(361));
    
    \AHB_Master_Out_pad[334]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(334));
    
    \AHB_Master_Out_pad[24]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[20]\, PAD => 
        AHB_Master_Out(24));
    
    \AHB_Master_In_pad[18]\ : INBUF
      port map(PAD => AHB_Master_In(18), Y => 
        \AHB_Master_In_c[18]\);
    
    \apbo_pad[35]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(35));
    
    \apbi_pad[51]\ : INBUF
      port map(PAD => apbi(51), Y => \apbi_c[51]\);
    
    \AHB_Master_Out_pad[253]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(253));
    
    \AHB_Master_Out_pad[177]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(177));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \apbo_pad[21]\ : OUTBUF
      port map(D => \apbo.prdata_c[21]\, PAD => apbo(21));
    
    \apbi_pad[55]\ : INBUF
      port map(PAD => apbi(55), Y => \apbi_c[55]\);
    
    \AHB_Master_Out_pad[151]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(151));
    
    \apbo_pad[25]\ : OUTBUF
      port map(D => \apbo.prdata_c[25]\, PAD => apbo(25));
    
    \apbo_pad[17]\ : OUTBUF
      port map(D => \apbo.prdata_c[17]\, PAD => apbo(17));
    
    \apbo_pad[120]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(120));
    
    \AHB_Master_Out_pad[300]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(300));
    
    data_shaping_BW_pad : OUTBUF
      port map(D => data_shaping_BW_c, PAD => data_shaping_BW);
    
    \apbi_pad[73]\ : INBUF
      port map(PAD => apbi(73), Y => \apbi_c[73]\);
    
    \AHB_Master_Out_pad[96]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(96));
    
    \AHB_Master_Out_pad[216]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(216));
    
    \apbo_pad[4]\ : OUTBUF
      port map(D => \apbo.prdata_c[4]\, PAD => apbo(4));
    
    \AHB_Master_Out_pad[226]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(226));
    
    \AHB_Master_Out_pad[42]\ : OUTBUF
      port map(D => \AHB_Master_Out.hburst_c[2]\, PAD => 
        AHB_Master_Out(42));
    
    \AHB_Master_Out_pad[246]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(246));
    
    \AHB_Master_Out_pad[260]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(260));
    
    \AHB_Master_Out_pad[118]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(118));
    
    \apbo_pad[61]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(61));
    
    \AHB_Master_Out_pad[294]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(294));
    
    \AHB_Master_Out_pad[165]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(165));
    
    \AHB_Master_Out_pad[128]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(128));
    
    \apbo_pad[65]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(65));
    
    \AHB_Master_Out_pad[148]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(148));
    
    \apbo_pad[13]\ : OUTBUF
      port map(D => \apbo.prdata_c[13]\, PAD => apbo(13));
    
    \AHB_Master_Out_pad[97]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(97));
    
    \apbi_pad[80]\ : INBUF
      port map(PAD => apbi(80), Y => \apbi_c[80]\);
    
    \AHB_Master_Out_pad[235]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(235));
    
    \apbo_pad[101]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(101));
    
    \AHB_Master_Out_pad[293]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(293));
    
    \AHB_Master_Out_pad[191]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(191));
    
    \AHB_Master_Out_pad[99]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(99));
    
    \apbo_pad[59]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(59));
    
    \apbo_pad[47]\ : OUTBUF
      port map(D => \apbo.pirq_c[15]\, PAD => apbo(47));
    
    \AHB_Master_Out_pad[266]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(266));
    
    \AHB_Master_Out_pad[23]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[19]\, PAD => 
        AHB_Master_Out(23));
    
    \apbo_pad[94]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(94));
    
    \apbo_pad[105]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(105));
    
    \AHB_Master_Out_pad[157]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(157));
    
    \AHB_Master_Out_pad[313]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(313));
    
    \AHB_Master_Out_pad[168]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(168));
    
    \AHB_Master_Out_pad[323]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(323));
    
    \AHB_Master_Out_pad[102]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(102));
    
    \AHB_Master_Out_pad[343]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(343));
    
    \apbo_pad[5]\ : OUTBUF
      port map(D => \apbo.prdata_c[5]\, PAD => apbo(5));
    
    \apbi_pad[81]\ : INBUF
      port map(PAD => apbi(81), Y => \apbi_c[81]\);
    
    \apbo_pad[43]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(43));
    
    lpp_top_apbreg_1 : lpp_top_apbreg
      port map(status_full_ack(3) => \status_full_ack[3]\, 
        status_full_ack(2) => \status_full_ack[2]\, 
        status_full_ack(1) => \status_full_ack[1]\, 
        status_full_ack(0) => \status_full_ack[0]\, prdata_c(31)
         => \apbo.prdata_c[31]\, prdata_c(30) => 
        \apbo.prdata_c[30]\, prdata_c(29) => \apbo.prdata_c[29]\, 
        prdata_c(28) => \apbo.prdata_c[28]\, prdata_c(27) => 
        \apbo.prdata_c[27]\, prdata_c(26) => \apbo.prdata_c[26]\, 
        prdata_c(25) => \apbo.prdata_c[25]\, prdata_c(24) => 
        \apbo.prdata_c[24]\, prdata_c(23) => \apbo.prdata_c[23]\, 
        prdata_c(22) => \apbo.prdata_c[22]\, prdata_c(21) => 
        \apbo.prdata_c[21]\, prdata_c(20) => \apbo.prdata_c[20]\, 
        prdata_c(19) => \apbo.prdata_c[19]\, prdata_c(18) => 
        \apbo.prdata_c[18]\, prdata_c(17) => \apbo.prdata_c[17]\, 
        prdata_c(16) => \apbo.prdata_c[16]\, prdata_c(15) => 
        \apbo.prdata_c[15]\, prdata_c(14) => \apbo.prdata_c[14]\, 
        prdata_c(13) => \apbo.prdata_c[13]\, prdata_c(12) => 
        \apbo.prdata_c[12]\, prdata_c(11) => \apbo.prdata_c[11]\, 
        prdata_c(10) => \apbo.prdata_c[10]\, prdata_c(9) => 
        \apbo.prdata_c[9]\, prdata_c(8) => \apbo.prdata_c[8]\, 
        prdata_c(7) => \apbo.prdata_c[7]\, prdata_c(6) => 
        \apbo.prdata_c[6]\, prdata_c(5) => \apbo.prdata_c[5]\, 
        prdata_c(4) => \apbo.prdata_c[4]\, prdata_c(3) => 
        \apbo.prdata_c[3]\, prdata_c(2) => \apbo.prdata_c[2]\, 
        prdata_c(1) => \apbo.prdata_c[1]\, prdata_c(0) => 
        \apbo.prdata_c[0]\, pirq_c(15) => \apbo.pirq_c[15]\, 
        addr_data_f2(31) => \addr_data_f2[31]\, addr_data_f2(30)
         => \addr_data_f2[30]\, addr_data_f2(29) => 
        \addr_data_f2[29]\, addr_data_f2(28) => 
        \addr_data_f2[28]\, addr_data_f2(27) => 
        \addr_data_f2[27]\, addr_data_f2(26) => 
        \addr_data_f2[26]\, addr_data_f2(25) => 
        \addr_data_f2[25]\, addr_data_f2(24) => 
        \addr_data_f2[24]\, addr_data_f2(23) => 
        \addr_data_f2[23]\, addr_data_f2(22) => 
        \addr_data_f2[22]\, addr_data_f2(21) => 
        \addr_data_f2[21]\, addr_data_f2(20) => 
        \addr_data_f2[20]\, addr_data_f2(19) => 
        \addr_data_f2[19]\, addr_data_f2(18) => 
        \addr_data_f2[18]\, addr_data_f2(17) => 
        \addr_data_f2[17]\, addr_data_f2(16) => 
        \addr_data_f2[16]\, addr_data_f2(15) => 
        \addr_data_f2[15]\, addr_data_f2(14) => 
        \addr_data_f2[14]\, addr_data_f2(13) => 
        \addr_data_f2[13]\, addr_data_f2(12) => 
        \addr_data_f2[12]\, addr_data_f2(11) => 
        \addr_data_f2[11]\, addr_data_f2(10) => 
        \addr_data_f2[10]\, addr_data_f2(9) => \addr_data_f2[9]\, 
        addr_data_f2(8) => \addr_data_f2[8]\, addr_data_f2(7) => 
        \addr_data_f2[7]\, addr_data_f2(6) => \addr_data_f2[6]\, 
        addr_data_f2(5) => \addr_data_f2[5]\, addr_data_f2(4) => 
        \addr_data_f2[4]\, addr_data_f2(3) => \addr_data_f2[3]\, 
        addr_data_f2(2) => \addr_data_f2[2]\, addr_data_f2(1) => 
        \addr_data_f2[1]\, addr_data_f2(0) => \addr_data_f2[0]\, 
        status_new_err_3 => \status_new_err[3]\, 
        status_new_err_0_2 => \status_new_err[2]\, 
        status_new_err_0_0 => \status_new_err[0]\, 
        status_new_err_0_1 => \status_new_err[1]\, 
        status_full_err_0(3) => \status_full_err[3]\, 
        status_full_err_0(2) => \status_full_err[2]\, 
        status_full_err_0(1) => \status_full_err[1]\, 
        status_full_err_0(0) => \status_full_err[0]\, 
        status_full(3) => \status_full[3]\, status_full(2) => 
        \status_full[2]\, status_full(1) => \status_full[1]\, 
        status_full(0) => \status_full[0]\, addr_data_f3(31) => 
        \addr_data_f3[31]\, addr_data_f3(30) => 
        \addr_data_f3[30]\, addr_data_f3(29) => 
        \addr_data_f3[29]\, addr_data_f3(28) => 
        \addr_data_f3[28]\, addr_data_f3(27) => 
        \addr_data_f3[27]\, addr_data_f3(26) => 
        \addr_data_f3[26]\, addr_data_f3(25) => 
        \addr_data_f3[25]\, addr_data_f3(24) => 
        \addr_data_f3[24]\, addr_data_f3(23) => 
        \addr_data_f3[23]\, addr_data_f3(22) => 
        \addr_data_f3[22]\, addr_data_f3(21) => 
        \addr_data_f3[21]\, addr_data_f3(20) => 
        \addr_data_f3[20]\, addr_data_f3(19) => 
        \addr_data_f3[19]\, addr_data_f3(18) => 
        \addr_data_f3[18]\, addr_data_f3(17) => 
        \addr_data_f3[17]\, addr_data_f3(16) => 
        \addr_data_f3[16]\, addr_data_f3(15) => 
        \addr_data_f3[15]\, addr_data_f3(14) => 
        \addr_data_f3[14]\, addr_data_f3(13) => 
        \addr_data_f3[13]\, addr_data_f3(12) => 
        \addr_data_f3[12]\, addr_data_f3(11) => 
        \addr_data_f3[11]\, addr_data_f3(10) => 
        \addr_data_f3[10]\, addr_data_f3(9) => \addr_data_f3[9]\, 
        addr_data_f3(8) => \addr_data_f3[8]\, addr_data_f3(7) => 
        \addr_data_f3[7]\, addr_data_f3(6) => \addr_data_f3[6]\, 
        addr_data_f3(5) => \addr_data_f3[5]\, addr_data_f3(4) => 
        \addr_data_f3[4]\, addr_data_f3(3) => \addr_data_f3[3]\, 
        addr_data_f3(2) => \addr_data_f3[2]\, addr_data_f3(1) => 
        \addr_data_f3[1]\, addr_data_f3(0) => \addr_data_f3[0]\, 
        nb_burst_available(10) => \nb_burst_available[10]\, 
        nb_burst_available(9) => \nb_burst_available[9]\, 
        nb_burst_available(8) => \nb_burst_available[8]\, 
        nb_burst_available(7) => \nb_burst_available[7]\, 
        nb_burst_available(6) => \nb_burst_available[6]\, 
        nb_burst_available(5) => \nb_burst_available[5]\, 
        nb_burst_available(4) => \nb_burst_available[4]\, 
        nb_burst_available(3) => \nb_burst_available[3]\, 
        nb_burst_available(2) => \nb_burst_available[2]\, 
        nb_burst_available(1) => \nb_burst_available[1]\, 
        nb_burst_available(0) => \nb_burst_available[0]\, 
        addr_data_f1(31) => \addr_data_f1[31]\, addr_data_f1(30)
         => \addr_data_f1[30]\, addr_data_f1(29) => 
        \addr_data_f1[29]\, addr_data_f1(28) => 
        \addr_data_f1[28]\, addr_data_f1(27) => 
        \addr_data_f1[27]\, addr_data_f1(26) => 
        \addr_data_f1[26]\, addr_data_f1(25) => 
        \addr_data_f1[25]\, addr_data_f1(24) => 
        \addr_data_f1[24]\, addr_data_f1(23) => 
        \addr_data_f1[23]\, addr_data_f1(22) => 
        \addr_data_f1[22]\, addr_data_f1(21) => 
        \addr_data_f1[21]\, addr_data_f1(20) => 
        \addr_data_f1[20]\, addr_data_f1(19) => 
        \addr_data_f1[19]\, addr_data_f1(18) => 
        \addr_data_f1[18]\, addr_data_f1(17) => 
        \addr_data_f1[17]\, addr_data_f1(16) => 
        \addr_data_f1[16]\, addr_data_f1(15) => 
        \addr_data_f1[15]\, addr_data_f1(14) => 
        \addr_data_f1[14]\, addr_data_f1(13) => 
        \addr_data_f1[13]\, addr_data_f1(12) => 
        \addr_data_f1[12]\, addr_data_f1(11) => 
        \addr_data_f1[11]\, addr_data_f1(10) => 
        \addr_data_f1[10]\, addr_data_f1(9) => \addr_data_f1[9]\, 
        addr_data_f1(8) => \addr_data_f1[8]\, addr_data_f1(7) => 
        \addr_data_f1[7]\, addr_data_f1(6) => \addr_data_f1[6]\, 
        addr_data_f1(5) => \addr_data_f1[5]\, addr_data_f1(4) => 
        \addr_data_f1[4]\, addr_data_f1(3) => \addr_data_f1[3]\, 
        addr_data_f1(2) => \addr_data_f1[2]\, addr_data_f1(1) => 
        \addr_data_f1[1]\, addr_data_f1(0) => \addr_data_f1[0]\, 
        delta_f2_f1(9) => \delta_f2_f1[9]\, delta_f2_f1(8) => 
        \delta_f2_f1[8]\, delta_f2_f1(7) => \delta_f2_f1[7]\, 
        delta_f2_f1(6) => \delta_f2_f1[6]\, delta_f2_f1(5) => 
        \delta_f2_f1[5]\, delta_f2_f1(4) => \delta_f2_f1[4]\, 
        delta_f2_f1(3) => \delta_f2_f1[3]\, delta_f2_f1(2) => 
        \delta_f2_f1[2]\, delta_f2_f1(1) => \delta_f2_f1[1]\, 
        delta_f2_f1(0) => \delta_f2_f1[0]\, addr_data_f0(31) => 
        \addr_data_f0[31]\, addr_data_f0(30) => 
        \addr_data_f0[30]\, addr_data_f0(29) => 
        \addr_data_f0[29]\, addr_data_f0(28) => 
        \addr_data_f0[28]\, addr_data_f0(27) => 
        \addr_data_f0[27]\, addr_data_f0(26) => 
        \addr_data_f0[26]\, addr_data_f0(25) => 
        \addr_data_f0[25]\, addr_data_f0(24) => 
        \addr_data_f0[24]\, addr_data_f0(23) => 
        \addr_data_f0[23]\, addr_data_f0(22) => 
        \addr_data_f0[22]\, addr_data_f0(21) => 
        \addr_data_f0[21]\, addr_data_f0(20) => 
        \addr_data_f0[20]\, addr_data_f0(19) => 
        \addr_data_f0[19]\, addr_data_f0(18) => 
        \addr_data_f0[18]\, addr_data_f0(17) => 
        \addr_data_f0[17]\, addr_data_f0(16) => 
        \addr_data_f0[16]\, addr_data_f0(15) => 
        \addr_data_f0[15]\, addr_data_f0(14) => 
        \addr_data_f0[14]\, addr_data_f0(13) => 
        \addr_data_f0[13]\, addr_data_f0(12) => 
        \addr_data_f0[12]\, addr_data_f0(11) => 
        \addr_data_f0[11]\, addr_data_f0(10) => 
        \addr_data_f0[10]\, addr_data_f0(9) => \addr_data_f0[9]\, 
        addr_data_f0(8) => \addr_data_f0[8]\, addr_data_f0(7) => 
        \addr_data_f0[7]\, addr_data_f0(6) => \addr_data_f0[6]\, 
        addr_data_f0(5) => \addr_data_f0[5]\, addr_data_f0(4) => 
        \addr_data_f0[4]\, addr_data_f0(3) => \addr_data_f0[3]\, 
        addr_data_f0(2) => \addr_data_f0[2]\, addr_data_f0(1) => 
        \addr_data_f0[1]\, addr_data_f0(0) => \addr_data_f0[0]\, 
        delta_f2_f0(9) => \delta_f2_f0[9]\, delta_f2_f0(8) => 
        \delta_f2_f0[8]\, delta_f2_f0(7) => \delta_f2_f0[7]\, 
        delta_f2_f0(6) => \delta_f2_f0[6]\, delta_f2_f0(5) => 
        \delta_f2_f0[5]\, delta_f2_f0(4) => \delta_f2_f0[4]\, 
        delta_f2_f0(3) => \delta_f2_f0[3]\, delta_f2_f0(2) => 
        \delta_f2_f0[2]\, delta_f2_f0(1) => \delta_f2_f0[1]\, 
        delta_f2_f0(0) => \delta_f2_f0[0]\, delta_snapshot(15)
         => \delta_snapshot[15]\, delta_snapshot(14) => 
        \delta_snapshot[14]\, delta_snapshot(13) => 
        \delta_snapshot[13]\, delta_snapshot(12) => 
        \delta_snapshot[12]\, delta_snapshot(11) => 
        \delta_snapshot[11]\, delta_snapshot(10) => 
        \delta_snapshot[10]\, delta_snapshot(9) => 
        \delta_snapshot[9]\, delta_snapshot(8) => 
        \delta_snapshot[8]\, delta_snapshot(7) => 
        \delta_snapshot[7]\, delta_snapshot(6) => 
        \delta_snapshot[6]\, delta_snapshot(5) => 
        \delta_snapshot[5]\, delta_snapshot(4) => 
        \delta_snapshot[4]\, delta_snapshot(3) => 
        \delta_snapshot[3]\, delta_snapshot(2) => 
        \delta_snapshot[2]\, delta_snapshot(1) => 
        \delta_snapshot[1]\, delta_snapshot(0) => 
        \delta_snapshot[0]\, nb_snapshot_param(10) => 
        \nb_snapshot_param[10]\, nb_snapshot_param(9) => 
        \nb_snapshot_param[9]\, nb_snapshot_param(8) => 
        \nb_snapshot_param[8]\, nb_snapshot_param(7) => 
        \nb_snapshot_param[7]\, nb_snapshot_param(6) => 
        \nb_snapshot_param[6]\, nb_snapshot_param(5) => 
        \nb_snapshot_param[5]\, nb_snapshot_param(4) => 
        \nb_snapshot_param[4]\, nb_snapshot_param(3) => 
        \nb_snapshot_param[3]\, nb_snapshot_param(2) => 
        \nb_snapshot_param[2]\, nb_snapshot_param(1) => 
        \nb_snapshot_param[1]\, nb_snapshot_param(0) => 
        \nb_snapshot_param[0]\, apbi_c_81 => \apbi_c[81]\, 
        apbi_c_80 => \apbi_c[80]\, apbi_c_79 => \apbi_c[79]\, 
        apbi_c_78 => \apbi_c[78]\, apbi_c_77 => \apbi_c[77]\, 
        apbi_c_76 => \apbi_c[76]\, apbi_c_75 => \apbi_c[75]\, 
        apbi_c_74 => \apbi_c[74]\, apbi_c_73 => \apbi_c[73]\, 
        apbi_c_72 => \apbi_c[72]\, apbi_c_71 => \apbi_c[71]\, 
        apbi_c_70 => \apbi_c[70]\, apbi_c_69 => \apbi_c[69]\, 
        apbi_c_68 => \apbi_c[68]\, apbi_c_67 => \apbi_c[67]\, 
        apbi_c_66 => \apbi_c[66]\, apbi_c_65 => \apbi_c[65]\, 
        apbi_c_64 => \apbi_c[64]\, apbi_c_63 => \apbi_c[63]\, 
        apbi_c_62 => \apbi_c[62]\, apbi_c_61 => \apbi_c[61]\, 
        apbi_c_60 => \apbi_c[60]\, apbi_c_59 => \apbi_c[59]\, 
        apbi_c_58 => \apbi_c[58]\, apbi_c_57 => \apbi_c[57]\, 
        apbi_c_56 => \apbi_c[56]\, apbi_c_55 => \apbi_c[55]\, 
        apbi_c_24 => \apbi_c[24]\, apbi_c_23 => \apbi_c[23]\, 
        apbi_c_0 => \apbi_c[0]\, apbi_c_50 => \apbi_c[50]\, 
        apbi_c_51 => \apbi_c[51]\, apbi_c_52 => \apbi_c[52]\, 
        apbi_c_16 => \apbi_c[16]\, apbi_c_49 => \apbi_c[49]\, 
        apbi_c_22 => \apbi_c[22]\, apbi_c_20 => \apbi_c[20]\, 
        apbi_c_19 => \apbi_c[19]\, apbi_c_21 => \apbi_c[21]\, 
        apbi_c_54 => \apbi_c[54]\, apbi_c_53 => \apbi_c[53]\, 
        data_shaping_R0 => data_shaping_R0, data_shaping_R1 => 
        data_shaping_R1, enable_f0 => enable_f0, 
        data_shaping_BW_c => data_shaping_BW_c, burst_f2 => 
        burst_f2, burst_f1 => burst_f1, burst_f0 => burst_f0, 
        enable_f3 => enable_f3, enable_f2 => enable_f2, 
        data_shaping_SP1 => data_shaping_SP1, enable_f1 => 
        enable_f1, data_shaping_SP0 => data_shaping_SP0, 
        data_shaping_R1_0 => data_shaping_R1_0, HRESETn_c => 
        HRESETn_c, HCLK_c => HCLK_c, data_shaping_R0_0 => 
        data_shaping_R0_0);
    
    \AHB_Master_Out_pad[78]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[31]\, PAD => 
        AHB_Master_Out(78));
    
    \AHB_Master_Out_pad[271]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(271));
    
    cnv_pad : OUTBUF
      port map(D => cnv_c, PAD => cnv);
    
    \AHB_Master_Out_pad[302]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(302));
    
    \AHB_Master_Out_pad[88]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(88));
    
    \AHB_Master_Out_pad[363]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(363));
    
    \AHB_Master_Out_pad[218]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(218));
    
    \AHB_Master_Out_pad[197]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(197));
    
    \apbo_pad[104]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(104));
    
    \AHB_Master_Out_pad[70]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[23]\, PAD => 
        AHB_Master_Out(70));
    
    \AHB_Master_Out_pad[228]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(228));
    
    \AHB_Master_Out_pad[248]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(248));
    
    \AHB_Master_Out_pad[285]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(285));
    
    \sdo_pad[3]\ : INBUF
      port map(PAD => sdo(3), Y => \sdo_c[3]\);
    
    \AHB_Master_Out_pad[80]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(80));
    
    \AHB_Master_Out_pad[309]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(309));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \apbo_pad[82]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(82));
    
    \apbi_pad[67]\ : INBUF
      port map(PAD => apbi(67), Y => \apbi_c[67]\);
    
    \AHB_Master_Out_pad[119]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(119));
    
    \apbo_pad[0]\ : OUTBUF
      port map(D => \apbo.prdata_c[0]\, PAD => apbo(0));
    
    \AHB_Master_Out_pad[129]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(129));
    
    \AHB_Master_Out_pad[149]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(149));
    
    \AHB_Master_Out_pad[58]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[11]\, PAD => 
        AHB_Master_Out(58));
    
    \AHB_Master_Out_pad[270]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(270));
    
    \AHB_Master_Out_pad[268]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(268));
    
    \AHB_Master_Out_pad[251]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(251));
    
    \AHB_Master_Out_pad[237]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(237));
    
    \AHB_Master_Out_pad[175]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(175));
    
    \AHB_Master_Out_pad[11]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[7]\, PAD => 
        AHB_Master_Out(11));
    
    \apbi_pad[63]\ : INBUF
      port map(PAD => apbi(63), Y => \apbi_c[63]\);
    
    \AHB_Master_Out_pad[76]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[29]\, PAD => 
        AHB_Master_Out(76));
    
    \AHB_Master_Out_pad[357]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(357));
    
    \apbo_pad[80]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(80));
    
    \AHB_Master_Out_pad[44]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(44));
    
    \AHB_Master_Out_pad[310]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(310));
    
    \AHB_Master_Out_pad[86]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(86));
    
    \AHB_Master_Out_pad[50]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[3]\, PAD => 
        AHB_Master_Out(50));
    
    \AHB_Master_Out_pad[320]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(320));
    
    \AHB_Master_Out_pad[239]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(239));
    
    \AHB_Master_Out_pad[202]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(202));
    
    \sdo_pad[5]\ : INBUF
      port map(PAD => sdo(5), Y => \sdo_c[5]\);
    
    lpp_top_lfr_wf_picker_ip_1 : lpp_top_lfr_wf_picker_ip
      port map(nb_snapshot_param(10) => \nb_snapshot_param[10]\, 
        nb_snapshot_param(9) => \nb_snapshot_param[9]\, 
        nb_snapshot_param(8) => \nb_snapshot_param[8]\, 
        nb_snapshot_param(7) => \nb_snapshot_param[7]\, 
        nb_snapshot_param(6) => \nb_snapshot_param[6]\, 
        nb_snapshot_param(5) => \nb_snapshot_param[5]\, 
        nb_snapshot_param(4) => \nb_snapshot_param[4]\, 
        nb_snapshot_param(3) => \nb_snapshot_param[3]\, 
        nb_snapshot_param(2) => \nb_snapshot_param[2]\, 
        nb_snapshot_param(1) => \nb_snapshot_param[1]\, 
        nb_snapshot_param(0) => \nb_snapshot_param[0]\, 
        delta_f2_f0(9) => \delta_f2_f0[9]\, delta_f2_f0(8) => 
        \delta_f2_f0[8]\, delta_f2_f0(7) => \delta_f2_f0[7]\, 
        delta_f2_f0(6) => \delta_f2_f0[6]\, delta_f2_f0(5) => 
        \delta_f2_f0[5]\, delta_f2_f0(4) => \delta_f2_f0[4]\, 
        delta_f2_f0(3) => \delta_f2_f0[3]\, delta_f2_f0(2) => 
        \delta_f2_f0[2]\, delta_f2_f0(1) => \delta_f2_f0[1]\, 
        delta_f2_f0(0) => \delta_f2_f0[0]\, delta_snapshot(15)
         => \delta_snapshot[15]\, delta_snapshot(14) => 
        \delta_snapshot[14]\, delta_snapshot(13) => 
        \delta_snapshot[13]\, delta_snapshot(12) => 
        \delta_snapshot[12]\, delta_snapshot(11) => 
        \delta_snapshot[11]\, delta_snapshot(10) => 
        \delta_snapshot[10]\, delta_snapshot(9) => 
        \delta_snapshot[9]\, delta_snapshot(8) => 
        \delta_snapshot[8]\, delta_snapshot(7) => 
        \delta_snapshot[7]\, delta_snapshot(6) => 
        \delta_snapshot[6]\, delta_snapshot(5) => 
        \delta_snapshot[5]\, delta_snapshot(4) => 
        \delta_snapshot[4]\, delta_snapshot(3) => 
        \delta_snapshot[3]\, delta_snapshot(2) => 
        \delta_snapshot[2]\, delta_snapshot(1) => 
        \delta_snapshot[1]\, delta_snapshot(0) => 
        \delta_snapshot[0]\, delta_f2_f1(9) => \delta_f2_f1[9]\, 
        delta_f2_f1(8) => \delta_f2_f1[8]\, delta_f2_f1(7) => 
        \delta_f2_f1[7]\, delta_f2_f1(6) => \delta_f2_f1[6]\, 
        delta_f2_f1(5) => \delta_f2_f1[5]\, delta_f2_f1(4) => 
        \delta_f2_f1[4]\, delta_f2_f1(3) => \delta_f2_f1[3]\, 
        delta_f2_f1(2) => \delta_f2_f1[2]\, delta_f2_f1(1) => 
        \delta_f2_f1[1]\, delta_f2_f1(0) => \delta_f2_f1[0]\, 
        status_new_err(3) => \status_new_err[3]\, 
        status_new_err(2) => \status_new_err[2]\, 
        status_new_err(1) => \status_new_err[1]\, 
        status_new_err(0) => \status_new_err[0]\, hwdata_c(31)
         => \AHB_Master_Out.hwdata_c[31]\, hwdata_c(30) => 
        \AHB_Master_Out.hwdata_c[30]\, hwdata_c(29) => 
        \AHB_Master_Out.hwdata_c[29]\, hwdata_c(28) => 
        \AHB_Master_Out.hwdata_c[28]\, hwdata_c(27) => 
        \AHB_Master_Out.hwdata_c[27]\, hwdata_c(26) => 
        \AHB_Master_Out.hwdata_c[26]\, hwdata_c(25) => 
        \AHB_Master_Out.hwdata_c[25]\, hwdata_c(24) => 
        \AHB_Master_Out.hwdata_c[24]\, hwdata_c(23) => 
        \AHB_Master_Out.hwdata_c[23]\, hwdata_c(22) => 
        \AHB_Master_Out.hwdata_c[22]\, hwdata_c(21) => 
        \AHB_Master_Out.hwdata_c[21]\, hwdata_c(20) => 
        \AHB_Master_Out.hwdata_c[20]\, hwdata_c(19) => 
        \AHB_Master_Out.hwdata_c[19]\, hwdata_c(18) => 
        \AHB_Master_Out.hwdata_c[18]\, hwdata_c(17) => 
        \AHB_Master_Out.hwdata_c[17]\, hwdata_c(16) => 
        \AHB_Master_Out.hwdata_c[16]\, hwdata_c(15) => 
        \AHB_Master_Out.hwdata_c[15]\, hwdata_c(14) => 
        \AHB_Master_Out.hwdata_c[14]\, hwdata_c(13) => 
        \AHB_Master_Out.hwdata_c[13]\, hwdata_c(12) => 
        \AHB_Master_Out.hwdata_c[12]\, hwdata_c(11) => 
        \AHB_Master_Out.hwdata_c[11]\, hwdata_c(10) => 
        \AHB_Master_Out.hwdata_c[10]\, hwdata_c(9) => 
        \AHB_Master_Out.hwdata_c[9]\, hwdata_c(8) => 
        \AHB_Master_Out.hwdata_c[8]\, hwdata_c(7) => 
        \AHB_Master_Out.hwdata_c[7]\, hwdata_c(6) => 
        \AHB_Master_Out.hwdata_c[6]\, hwdata_c(5) => 
        \AHB_Master_Out.hwdata_c[5]\, hwdata_c(4) => 
        \AHB_Master_Out.hwdata_c[4]\, hwdata_c(3) => 
        \AHB_Master_Out.hwdata_c[3]\, hwdata_c(2) => 
        \AHB_Master_Out.hwdata_c[2]\, hwdata_c(1) => 
        \AHB_Master_Out.hwdata_c[1]\, hwdata_c(0) => 
        \AHB_Master_Out.hwdata_c[0]\, addr_data_f0(31) => 
        \addr_data_f0[31]\, addr_data_f0(30) => 
        \addr_data_f0[30]\, addr_data_f0(29) => 
        \addr_data_f0[29]\, addr_data_f0(28) => 
        \addr_data_f0[28]\, addr_data_f0(27) => 
        \addr_data_f0[27]\, addr_data_f0(26) => 
        \addr_data_f0[26]\, addr_data_f0(25) => 
        \addr_data_f0[25]\, addr_data_f0(24) => 
        \addr_data_f0[24]\, addr_data_f0(23) => 
        \addr_data_f0[23]\, addr_data_f0(22) => 
        \addr_data_f0[22]\, addr_data_f0(21) => 
        \addr_data_f0[21]\, addr_data_f0(20) => 
        \addr_data_f0[20]\, addr_data_f0(19) => 
        \addr_data_f0[19]\, addr_data_f0(18) => 
        \addr_data_f0[18]\, addr_data_f0(17) => 
        \addr_data_f0[17]\, addr_data_f0(16) => 
        \addr_data_f0[16]\, addr_data_f0(15) => 
        \addr_data_f0[15]\, addr_data_f0(14) => 
        \addr_data_f0[14]\, addr_data_f0(13) => 
        \addr_data_f0[13]\, addr_data_f0(12) => 
        \addr_data_f0[12]\, addr_data_f0(11) => 
        \addr_data_f0[11]\, addr_data_f0(10) => 
        \addr_data_f0[10]\, addr_data_f0(9) => \addr_data_f0[9]\, 
        addr_data_f0(8) => \addr_data_f0[8]\, addr_data_f0(7) => 
        \addr_data_f0[7]\, addr_data_f0(6) => \addr_data_f0[6]\, 
        addr_data_f0(5) => \addr_data_f0[5]\, addr_data_f0(4) => 
        \addr_data_f0[4]\, addr_data_f0(3) => \addr_data_f0[3]\, 
        addr_data_f0(2) => \addr_data_f0[2]\, addr_data_f0(1) => 
        \addr_data_f0[1]\, addr_data_f0(0) => \addr_data_f0[0]\, 
        addr_data_f1(31) => \addr_data_f1[31]\, addr_data_f1(30)
         => \addr_data_f1[30]\, addr_data_f1(29) => 
        \addr_data_f1[29]\, addr_data_f1(28) => 
        \addr_data_f1[28]\, addr_data_f1(27) => 
        \addr_data_f1[27]\, addr_data_f1(26) => 
        \addr_data_f1[26]\, addr_data_f1(25) => 
        \addr_data_f1[25]\, addr_data_f1(24) => 
        \addr_data_f1[24]\, addr_data_f1(23) => 
        \addr_data_f1[23]\, addr_data_f1(22) => 
        \addr_data_f1[22]\, addr_data_f1(21) => 
        \addr_data_f1[21]\, addr_data_f1(20) => 
        \addr_data_f1[20]\, addr_data_f1(19) => 
        \addr_data_f1[19]\, addr_data_f1(18) => 
        \addr_data_f1[18]\, addr_data_f1(17) => 
        \addr_data_f1[17]\, addr_data_f1(16) => 
        \addr_data_f1[16]\, addr_data_f1(15) => 
        \addr_data_f1[15]\, addr_data_f1(14) => 
        \addr_data_f1[14]\, addr_data_f1(13) => 
        \addr_data_f1[13]\, addr_data_f1(12) => 
        \addr_data_f1[12]\, addr_data_f1(11) => 
        \addr_data_f1[11]\, addr_data_f1(10) => 
        \addr_data_f1[10]\, addr_data_f1(9) => \addr_data_f1[9]\, 
        addr_data_f1(8) => \addr_data_f1[8]\, addr_data_f1(7) => 
        \addr_data_f1[7]\, addr_data_f1(6) => \addr_data_f1[6]\, 
        addr_data_f1(5) => \addr_data_f1[5]\, addr_data_f1(4) => 
        \addr_data_f1[4]\, addr_data_f1(3) => \addr_data_f1[3]\, 
        addr_data_f1(2) => \addr_data_f1[2]\, addr_data_f1(1) => 
        \addr_data_f1[1]\, addr_data_f1(0) => \addr_data_f1[0]\, 
        addr_data_f2(31) => \addr_data_f2[31]\, addr_data_f2(30)
         => \addr_data_f2[30]\, addr_data_f2(29) => 
        \addr_data_f2[29]\, addr_data_f2(28) => 
        \addr_data_f2[28]\, addr_data_f2(27) => 
        \addr_data_f2[27]\, addr_data_f2(26) => 
        \addr_data_f2[26]\, addr_data_f2(25) => 
        \addr_data_f2[25]\, addr_data_f2(24) => 
        \addr_data_f2[24]\, addr_data_f2(23) => 
        \addr_data_f2[23]\, addr_data_f2(22) => 
        \addr_data_f2[22]\, addr_data_f2(21) => 
        \addr_data_f2[21]\, addr_data_f2(20) => 
        \addr_data_f2[20]\, addr_data_f2(19) => 
        \addr_data_f2[19]\, addr_data_f2(18) => 
        \addr_data_f2[18]\, addr_data_f2(17) => 
        \addr_data_f2[17]\, addr_data_f2(16) => 
        \addr_data_f2[16]\, addr_data_f2(15) => 
        \addr_data_f2[15]\, addr_data_f2(14) => 
        \addr_data_f2[14]\, addr_data_f2(13) => 
        \addr_data_f2[13]\, addr_data_f2(12) => 
        \addr_data_f2[12]\, addr_data_f2(11) => 
        \addr_data_f2[11]\, addr_data_f2(10) => 
        \addr_data_f2[10]\, addr_data_f2(9) => \addr_data_f2[9]\, 
        addr_data_f2(8) => \addr_data_f2[8]\, addr_data_f2(7) => 
        \addr_data_f2[7]\, addr_data_f2(6) => \addr_data_f2[6]\, 
        addr_data_f2(5) => \addr_data_f2[5]\, addr_data_f2(4) => 
        \addr_data_f2[4]\, addr_data_f2(3) => \addr_data_f2[3]\, 
        addr_data_f2(2) => \addr_data_f2[2]\, addr_data_f2(1) => 
        \addr_data_f2[1]\, addr_data_f2(0) => \addr_data_f2[0]\, 
        addr_data_f3(31) => \addr_data_f3[31]\, addr_data_f3(30)
         => \addr_data_f3[30]\, addr_data_f3(29) => 
        \addr_data_f3[29]\, addr_data_f3(28) => 
        \addr_data_f3[28]\, addr_data_f3(27) => 
        \addr_data_f3[27]\, addr_data_f3(26) => 
        \addr_data_f3[26]\, addr_data_f3(25) => 
        \addr_data_f3[25]\, addr_data_f3(24) => 
        \addr_data_f3[24]\, addr_data_f3(23) => 
        \addr_data_f3[23]\, addr_data_f3(22) => 
        \addr_data_f3[22]\, addr_data_f3(21) => 
        \addr_data_f3[21]\, addr_data_f3(20) => 
        \addr_data_f3[20]\, addr_data_f3(19) => 
        \addr_data_f3[19]\, addr_data_f3(18) => 
        \addr_data_f3[18]\, addr_data_f3(17) => 
        \addr_data_f3[17]\, addr_data_f3(16) => 
        \addr_data_f3[16]\, addr_data_f3(15) => 
        \addr_data_f3[15]\, addr_data_f3(14) => 
        \addr_data_f3[14]\, addr_data_f3(13) => 
        \addr_data_f3[13]\, addr_data_f3(12) => 
        \addr_data_f3[12]\, addr_data_f3(11) => 
        \addr_data_f3[11]\, addr_data_f3(10) => 
        \addr_data_f3[10]\, addr_data_f3(9) => \addr_data_f3[9]\, 
        addr_data_f3(8) => \addr_data_f3[8]\, addr_data_f3(7) => 
        \addr_data_f3[7]\, addr_data_f3(6) => \addr_data_f3[6]\, 
        addr_data_f3(5) => \addr_data_f3[5]\, addr_data_f3(4) => 
        \addr_data_f3[4]\, addr_data_f3(3) => \addr_data_f3[3]\, 
        addr_data_f3(2) => \addr_data_f3[2]\, addr_data_f3(1) => 
        \addr_data_f3[1]\, addr_data_f3(0) => \addr_data_f3[0]\, 
        status_full(3) => \status_full[3]\, status_full(2) => 
        \status_full[2]\, status_full(1) => \status_full[1]\, 
        status_full(0) => \status_full[0]\, status_full_err(3)
         => \status_full_err[3]\, status_full_err(2) => 
        \status_full_err[2]\, status_full_err(1) => 
        \status_full_err[1]\, status_full_err(0) => 
        \status_full_err[0]\, nb_burst_available(10) => 
        \nb_burst_available[10]\, nb_burst_available(9) => 
        \nb_burst_available[9]\, nb_burst_available(8) => 
        \nb_burst_available[8]\, nb_burst_available(7) => 
        \nb_burst_available[7]\, nb_burst_available(6) => 
        \nb_burst_available[6]\, nb_burst_available(5) => 
        \nb_burst_available[5]\, nb_burst_available(4) => 
        \nb_burst_available[4]\, nb_burst_available(3) => 
        \nb_burst_available[3]\, nb_burst_available(2) => 
        \nb_burst_available[2]\, nb_burst_available(1) => 
        \nb_burst_available[1]\, nb_burst_available(0) => 
        \nb_burst_available[0]\, haddr_c(31) => 
        \AHB_Master_Out.haddr_c[31]\, haddr_c(30) => 
        \AHB_Master_Out.haddr_c[30]\, haddr_c(29) => 
        \AHB_Master_Out.haddr_c[29]\, haddr_c(28) => 
        \AHB_Master_Out.haddr_c[28]\, haddr_c(27) => 
        \AHB_Master_Out.haddr_c[27]\, haddr_c(26) => 
        \AHB_Master_Out.haddr_c[26]\, haddr_c(25) => 
        \AHB_Master_Out.haddr_c[25]\, haddr_c(24) => 
        \AHB_Master_Out.haddr_c[24]\, haddr_c(23) => 
        \AHB_Master_Out.haddr_c[23]\, haddr_c(22) => 
        \AHB_Master_Out.haddr_c[22]\, haddr_c(21) => 
        \AHB_Master_Out.haddr_c[21]\, haddr_c(20) => 
        \AHB_Master_Out.haddr_c[20]\, haddr_c(19) => 
        \AHB_Master_Out.haddr_c[19]\, haddr_c(18) => 
        \AHB_Master_Out.haddr_c[18]\, haddr_c(17) => 
        \AHB_Master_Out.haddr_c[17]\, haddr_c(16) => 
        \AHB_Master_Out.haddr_c[16]\, haddr_c(15) => 
        \AHB_Master_Out.haddr_c[15]\, haddr_c(14) => 
        \AHB_Master_Out.haddr_c[14]\, haddr_c(13) => 
        \AHB_Master_Out.haddr_c[13]\, haddr_c(12) => 
        \AHB_Master_Out.haddr_c[12]\, haddr_c(11) => 
        \AHB_Master_Out.haddr_c[11]\, haddr_c(10) => 
        \AHB_Master_Out.haddr_c[10]\, haddr_c(9) => 
        \AHB_Master_Out.haddr_c[9]\, haddr_c(8) => 
        \AHB_Master_Out.haddr_c[8]\, haddr_c(7) => 
        \AHB_Master_Out.haddr_c[7]\, haddr_c(6) => 
        \AHB_Master_Out.haddr_c[6]\, haddr_c(5) => 
        \AHB_Master_Out.haddr_c[5]\, haddr_c(4) => 
        \AHB_Master_Out.haddr_c[4]\, haddr_c(3) => 
        \AHB_Master_Out.haddr_c[3]\, haddr_c(2) => 
        \AHB_Master_Out.haddr_c[2]\, haddr_c(1) => 
        \AHB_Master_Out.haddr_c[1]\, haddr_c(0) => 
        \AHB_Master_Out.haddr_c[0]\, AHB_Master_In_c_3 => 
        \AHB_Master_In_c[16]\, AHB_Master_In_c_0 => 
        \AHB_Master_In_c[13]\, AHB_Master_In_c_4 => 
        \AHB_Master_In_c[17]\, AHB_Master_In_c_5 => 
        \AHB_Master_In_c[18]\, hsize_c(1) => 
        \AHB_Master_Out.hsize_c[1]\, hsize_c(0) => 
        \AHB_Master_Out.hsize_c[0]\, htrans_c(1) => 
        \AHB_Master_Out.htrans_c[1]\, htrans_c(0) => 
        \AHB_Master_Out.htrans_c[0]\, hburst_c(2) => 
        \AHB_Master_Out.hburst_c[2]\, hburst_c(1) => 
        \AHB_Master_Out.hburst_c[1]\, hburst_c(0) => 
        \AHB_Master_Out.hburst_c[0]\, status_full_ack(3) => 
        \status_full_ack[3]\, status_full_ack(2) => 
        \status_full_ack[2]\, status_full_ack(1) => 
        \status_full_ack[1]\, status_full_ack(0) => 
        \status_full_ack[0]\, sdo_c(7) => \sdo_c[7]\, sdo_c(6)
         => \sdo_c[6]\, sdo_c(5) => \sdo_c[5]\, sdo_c(4) => 
        \sdo_c[4]\, sdo_c(3) => \sdo_c[3]\, sdo_c(2) => 
        \sdo_c[2]\, sdo_c(1) => \sdo_c[1]\, sdo_c(0) => 
        \sdo_c[0]\, coarse_time_0_c => coarse_time_0_c, enable_f0
         => enable_f0, data_shaping_R0 => data_shaping_R0, 
        data_shaping_R0_0 => data_shaping_R0_0, burst_f0 => 
        burst_f0, data_shaping_R1 => data_shaping_R1, 
        data_shaping_R1_0 => data_shaping_R1_0, enable_f1 => 
        enable_f1, burst_f1 => burst_f1, enable_f2 => enable_f2, 
        burst_f2 => burst_f2, enable_f3 => enable_f3, N_43 => 
        \lpp_top_lfr_wf_picker_ip_1.lpp_waveform_1.pp_waveform_dma_1.DMA2AHB_1.N_43\, 
        IdlePhase_RNI03G71 => IdlePhase_RNI03G71, hwrite_c => 
        \AHB_Master_Out.hwrite_c\, lpp_top_lfr_wf_picker_ip_GND
         => \GND\, lpp_top_lfr_wf_picker_ip_VCC => \VCC\, 
        cnv_run_c => cnv_run_c, sck_c => sck_c, cnv_c => cnv_c, 
        cnv_clk_c => cnv_clk_c, cnv_rstn_c => cnv_rstn_c, 
        data_shaping_SP0 => data_shaping_SP0, data_shaping_SP1
         => data_shaping_SP1, HRESETn_c => HRESETn_c, HCLK_c => 
        HCLK_c);
    
    \apbo_pad[38]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(38));
    
    \AHB_Master_Out_pad[340]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(340));
    
    \AHB_Master_Out_pad[169]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(169));
    
    \apbi_pad[58]\ : INBUF
      port map(PAD => apbi(58), Y => \apbi_c[58]\);
    
    \AHB_Master_Out_pad[77]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[30]\, PAD => 
        AHB_Master_Out(77));
    
    \apbo_pad[28]\ : OUTBUF
      port map(D => \apbo.prdata_c[28]\, PAD => apbo(28));
    
    \AHB_Master_Out_pad[104]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(104));
    
    \AHB_Master_Out_pad[351]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(351));
    
    \AHB_Master_Out_pad[276]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(276));
    
    \apbo_pad[118]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(118));
    
    \AHB_Master_Out_pad[87]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(87));
    
    \AHB_Master_Out_pad[79]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(79));
    
    \AHB_Master_Out_pad[178]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(178));
    
    \AHB_Master_Out_pad[130]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(130));
    
    \apbo_pad[81]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(81));
    
    \AHB_Master_Out_pad[291]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(291));
    
    \apbo_pad[85]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(85));
    
    \apbo_pad[97]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(97));
    
    \apbo_pad[68]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(68));
    
    \AHB_Master_Out_pad[89]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(89));
    
    \AHB_Master_Out_pad[360]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(360));
    
    \AHB_Master_Out_pad[305]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(305));
    
    \AHB_Master_Out_pad[136]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(136));
    
    \AHB_Master_Out_pad[56]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[9]\, PAD => 
        AHB_Master_Out(56));
    
    \apbo_pad[130]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(130));
    
    \AHB_Master_Out_pad[250]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(250));
    
    \apbo_pad[1]\ : OUTBUF
      port map(D => \apbo.prdata_c[1]\, PAD => apbo(1));
    
    \AHB_Master_Out_pad[155]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(155));
    
    \apbo_pad[8]\ : OUTBUF
      port map(D => \apbo.prdata_c[8]\, PAD => apbo(8));
    
    \AHB_Master_Out_pad[112]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(112));
    
    \AHB_Master_Out_pad[43]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(43));
    
    \AHB_Master_Out_pad[122]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(122));
    
    \apbo_pad[93]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(93));
    
    \AHB_Master_Out_pad[57]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[10]\, PAD => 
        AHB_Master_Out(57));
    
    \AHB_Master_Out_pad[287]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(287));
    
    \AHB_Master_Out_pad[142]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(142));
    
    \apbo_pad[123]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(123));
    
    \AHB_Master_Out_pad[59]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[12]\, PAD => 
        AHB_Master_Out(59));
    
    \AHB_Master_Out_pad[289]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(289));
    
    \AHB_Master_Out_pad[256]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(256));
    
    \AHB_Master_Out_pad[95]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(95));
    
    \AHB_Master_Out_pad[312]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(312));
    
    \apbo_pad[107]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(107));
    
    \AHB_Master_Out_pad[322]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(322));
    
    \AHB_Master_Out_pad[158]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(158));
    
    \AHB_Master_Out_pad[342]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(342));
    
    \AHB_Master_Out_pad[290]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(290));
    
    \AHB_Master_Out_pad[103]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(103));
    
    \apbo_pad[36]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(36));
    
    \apbi_pad[16]\ : INBUF
      port map(PAD => apbi(16), Y => \apbi_c[16]\);
    
    \AHB_Master_Out_pad[68]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[21]\, PAD => 
        AHB_Master_Out(68));
    
    \AHB_Master_Out_pad[195]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(195));
    
    \AHB_Master_Out_pad[21]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[17]\, PAD => 
        AHB_Master_Out(21));
    
    \apbi_pad[56]\ : INBUF
      port map(PAD => apbi(56), Y => \apbi_c[56]\);
    
    \AHB_Master_Out_pad[162]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(162));
    
    \apbo_pad[72]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(72));
    
    \apbo_pad[26]\ : OUTBUF
      port map(D => \apbo.prdata_c[26]\, PAD => apbo(26));
    
    \apbi_pad[79]\ : INBUF
      port map(PAD => apbi(79), Y => \apbi_c[79]\);
    
    \AHB_Master_Out_pad[180]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(180));
    
    \AHB_Master_Out_pad[278]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(278));
    
    \AHB_Master_Out_pad[319]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(319));
    
    \AHB_Master_Out_pad[329]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(329));
    
    \apbo_pad[111]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(111));
    
    \AHB_Master_Out_pad[60]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[13]\, PAD => 
        AHB_Master_Out(60));
    
    \AHB_Master_Out_pad[349]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(349));
    
    \AHB_Master_Out_pad[186]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(186));
    
    \apbo_pad[19]\ : OUTBUF
      port map(D => \apbo.prdata_c[19]\, PAD => apbo(19));
    
    \AHB_Master_Out_pad[92]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(92));
    
    \AHB_Master_Out_pad[296]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(296));
    
    \apbo_pad[66]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(66));
    
    \AHB_Master_Out_pad[362]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(362));
    
    \AHB_Master_Out_pad[353]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(353));
    
    \AHB_Master_Out_pad[306]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(306));
    
    \AHB_Master_Out_pad[179]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(179));
    
    \apbo_pad[70]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(70));
    
    \apbi_pad[22]\ : INBUF
      port map(PAD => apbi(22), Y => \apbi_c[22]\);
    
    \AHB_Master_Out_pad[198]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(198));
    
    \apbo_pad[115]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(115));
    
    \AHB_Master_Out_pad[38]\ : OUTBUF
      port map(D => \AHB_Master_Out.hsize_c[1]\, PAD => 
        AHB_Master_Out(38));
    
    \AHB_Master_Out_pad[369]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(369));
    
    \AHB_Master_Out_pad[212]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(212));
    
    \AHB_Master_Out_pad[222]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(222));
    
    \AHB_Master_Out_pad[66]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[19]\, PAD => 
        AHB_Master_Out(66));
    
    \AHB_Master_Out_pad[242]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(242));
    
    \apbi_pad[20]\ : INBUF
      port map(PAD => apbi(20), Y => \apbi_c[20]\);
    
    \AHB_Master_Out_pad[370]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(370));
    
    \apbo_pad[34]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(34));
    
    \AHB_Master_Out_pad[114]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(114));
    
    \apbo_pad[49]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(49));
    
    \AHB_Master_Out_pad[124]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(124));
    
    \apbo_pad[71]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(71));
    
    \apbi_pad[54]\ : INBUF
      port map(PAD => apbi(54), Y => \apbi_c[54]\);
    
    \AHB_Master_Out_pad[30]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[26]\, PAD => 
        AHB_Master_Out(30));
    
    \AHB_Master_Out_pad[258]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(258));
    
    \AHB_Master_Out_pad[144]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(144));
    
    \apbo_pad[75]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(75));
    
    \apbo_pad[24]\ : OUTBUF
      port map(D => \apbo.prdata_c[24]\, PAD => apbo(24));
    
    \AHB_Master_Out_pad[67]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[20]\, PAD => 
        AHB_Master_Out(67));
    
    \apbo_pad[114]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(114));
    
    \AHB_Master_Out_pad[304]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(304));
    
    \apbo_pad[3]\ : OUTBUF
      port map(D => \apbo.prdata_c[3]\, PAD => apbo(3));
    
    \AHB_Master_Out_pad[315]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(315));
    
    \AHB_Master_Out_pad[159]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(159));
    
    \AHB_Master_Out_pad[69]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[22]\, PAD => 
        AHB_Master_Out(69));
    
    \AHB_Master_Out_pad[325]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(325));
    
    \AHB_Master_Out_pad[262]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(262));
    
    \apbo_pad[64]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(64));
    
    \AHB_Master_Out_pad[345]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(345));
    
    \apbi_pad[21]\ : INBUF
      port map(PAD => apbi(21), Y => \apbi_c[21]\);
    
    \apbo_pad[88]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(88));
    
    \AHB_Master_Out_pad[164]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(164));
    
    \apbo_pad[2]\ : OUTBUF
      port map(D => \apbo.prdata_c[2]\, PAD => apbo(2));
    
    \AHB_Master_Out_pad[36]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwrite_c\, PAD => 
        AHB_Master_Out(36));
    
    \AHB_Master_Out_pad[338]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(338));
    
    \AHB_Master_Out_pad[298]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(298));
    
    \AHB_Master_Out_pad[75]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[28]\, PAD => 
        AHB_Master_Out(75));
    
    \AHB_Master_Out_pad[172]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(172));
    
    \AHB_Master_Out_pad[350]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(350));
    
    \apbo_pad[100]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(100));
    
    \AHB_Master_Out_pad[85]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(85));
    
    \AHB_Master_Out_pad[205]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(205));
    
    \sdo_pad[7]\ : INBUF
      port map(PAD => sdo(7), Y => \sdo_c[7]\);
    
    \apbo_pad[52]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(52));
    
    \AHB_Master_Out_pad[37]\ : OUTBUF
      port map(D => \AHB_Master_Out.hsize_c[0]\, PAD => 
        AHB_Master_Out(37));
    
    \AHB_Master_Out_pad[365]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(365));
    
    \AHB_Master_Out_pad[199]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(199));
    
    \apbi_pad[69]\ : INBUF
      port map(PAD => apbi(69), Y => \apbi_c[69]\);
    
    \AHB_Master_Out_pad[113]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(113));
    
    \AHB_Master_Out_pad[234]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(234));
    
    \AHB_Master_Out_pad[123]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(123));
    
    \apbo_pad[129]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(129));
    
    \AHB_Master_Out_pad[39]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(39));
    
    \AHB_Master_Out_pad[143]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(143));
    
    HRESETn_pad : CLKBUF
      port map(PAD => HRESETn, Y => HRESETn_c);
    
    \AHB_Master_Out_pad[94]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(94));
    
    \AHB_Master_Out_pad[72]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[25]\, PAD => 
        AHB_Master_Out(72));
    
    \AHB_Master_Out_pad[41]\ : OUTBUF
      port map(D => \AHB_Master_Out.hburst_c[1]\, PAD => 
        AHB_Master_Out(41));
    
    \apbo_pad[50]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(50));
    
    \AHB_Master_Out_pad[233]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(233));
    
    \AHB_Master_Out_pad[131]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(131));
    
    \AHB_Master_Out_pad[8]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[4]\, PAD => 
        AHB_Master_Out(8));
    
    \AHB_Master_Out_pad[82]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(82));
    
    \AHB_Master_Out_pad[55]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[8]\, PAD => 
        AHB_Master_Out(55));
    
    \AHB_Master_Out_pad[316]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(316));
    
    \AHB_Master_Out_pad[326]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(326));
    
    \AHB_Master_Out_pad[163]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(163));
    
    \AHB_Master_Out_pad[152]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(152));
    
    \AHB_Master_Out_pad[346]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(346));
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \apbo_pad[86]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(86));
    
    \sdo_pad[0]\ : INBUF
      port map(PAD => sdo(0), Y => \sdo_c[0]\);
    
    \apbo_pad[51]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(51));
    
    \apbo_pad[37]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(37));
    
    \apbo_pad[55]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(55));
    
    \apbi_pad[57]\ : INBUF
      port map(PAD => apbi(57), Y => \apbi_c[57]\);
    
    \apbo_pad[27]\ : OUTBUF
      port map(D => \apbo.prdata_c[27]\, PAD => apbo(27));
    
    \AHB_Master_Out_pad[52]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[5]\, PAD => 
        AHB_Master_Out(52));
    
    \AHB_Master_Out_pad[352]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(352));
    
    \apbo_pad[99]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(99));
    
    \apbo_pad[126]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(126));
    
    \AHB_Master_Out_pad[272]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(272));
    
    \AHB_Master_Out_pad[93]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(93));
    
    \AHB_Master_Out_pad[366]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(366));
    
    \AHB_Master_Out_pad[284]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(284));
    
    \apbo_pad[117]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(117));
    
    \AHB_Master_Out_pad[137]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(137));
    
    \apbo_pad[33]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(33));
    
    \AHB_Master_Out_pad[192]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(192));
    
    \AHB_Master_Out_pad[174]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(174));
    
    \apbo_pad[122]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(122));
    
    \apbo_pad[67]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(67));
    
    \apbi_pad[53]\ : INBUF
      port map(PAD => apbi(53), Y => \apbi_c[53]\);
    
    \apbo_pad[23]\ : OUTBUF
      port map(D => \apbo.prdata_c[23]\, PAD => apbo(23));
    
    \AHB_Master_Out_pad[359]\ : OUTBUF
      port map(D => \VCC\, PAD => AHB_Master_Out(359));
    
    \AHB_Master_Out_pad[314]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(314));
    
    \AHB_Master_Out_pad[324]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(324));
    
    \AHB_Master_Out_pad[283]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(283));
    
    \AHB_Master_Out_pad[207]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(207));
    
    \apbo_pad[78]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(78));
    
    \AHB_Master_Out_pad[344]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(344));
    
    \AHB_Master_Out_pad[181]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(181));
    
    \AHB_Master_Out_pad[209]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(209));
    
    \apbo_pad[63]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(63));
    
    \apbo_pad[84]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(84));
    
    \AHB_Master_Out_pad[364]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(364));
    
    \AHB_Master_Out_pad[252]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(252));
    
    \AHB_Master_Out_pad[100]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(100));
    
    \AHB_Master_Out_pad[215]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(215));
    
    \AHB_Master_Out_pad[225]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(225));
    
    \AHB_Master_Out_pad[65]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[18]\, PAD => 
        AHB_Master_Out(65));
    
    \AHB_Master_Out_pad[245]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(245));
    
    \apbi_pad[0]\ : INBUF
      port map(PAD => apbi(0), Y => \apbi_c[0]\);
    
    \AHB_Master_Out_pad[154]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(154));
    
    \AHB_Master_Out_pad[74]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[27]\, PAD => 
        AHB_Master_Out(74));
    
    \AHB_Master_Out_pad[106]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(106));
    
    \AHB_Master_Out_pad[187]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(187));
    
    \AHB_Master_Out_pad[84]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(84));
    
    \AHB_Master_Out_pad[173]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(173));
    
    \AHB_Master_Out_pad[18]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[14]\, PAD => 
        AHB_Master_Out(18));
    
    \AHB_Master_Out_pad[231]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(231));
    
    \AHB_Master_Out_pad[337]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(337));
    
    \AHB_Master_Out_pad[355]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(355));
    
    \AHB_Master_Out_pad[292]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(292));
    
    \AHB_Master_Out_pad[265]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(265));
    
    \AHB_Master_Out_pad[62]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[15]\, PAD => 
        AHB_Master_Out(62));
    
    \apbo_pad[76]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(76));
    
    \AHB_Master_Out_pad[10]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[6]\, PAD => 
        AHB_Master_Out(10));
    
    \AHB_Master_Out_pad[9]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[5]\, PAD => 
        AHB_Master_Out(9));
    
    \AHB_Master_Out_pad[194]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(194));
    
    \AHB_Master_Out_pad[35]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[31]\, PAD => 
        AHB_Master_Out(35));
    
    \AHB_Master_Out_pad[331]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(331));
    
    \apbi_pad[72]\ : INBUF
      port map(PAD => apbi(72), Y => \apbi_c[72]\);
    
    cnv_rstn_pad : INBUF
      port map(PAD => cnv_rstn, Y => cnv_rstn_c);
    
    \AHB_Master_Out_pad[54]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[7]\, PAD => 
        AHB_Master_Out(54));
    
    \apbo_pad[103]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(103));
    
    \AHB_Master_Out_pad[73]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[26]\, PAD => 
        AHB_Master_Out(73));
    
    \apbo_pad[9]\ : OUTBUF
      port map(D => \apbo.prdata_c[9]\, PAD => apbo(9));
    
    \apbo_pad[12]\ : OUTBUF
      port map(D => \apbo.prdata_c[12]\, PAD => apbo(12));
    
    \apbo_pad[110]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(110));
    
    \AHB_Master_Out_pad[153]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(153));
    
    \AHB_Master_Out_pad[83]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(83));
    
    \AHB_Master_Out_pad[5]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[1]\, PAD => 
        AHB_Master_Out(5));
    
    \AHB_Master_Out_pad[230]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(230));
    
    \apbo_pad[58]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(58));
    
    \apbi_pad[70]\ : INBUF
      port map(PAD => apbi(70), Y => \apbi_c[70]\);
    
    \AHB_Master_Out_pad[16]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[12]\, PAD => 
        AHB_Master_Out(16));
    
    \AHB_Master_Out_pad[135]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(135));
    
    \AHB_Master_Out_pad[32]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[28]\, PAD => 
        AHB_Master_Out(32));
    
    \AHB_Master_Out_pad[281]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(281));
    
    \apbo_pad[10]\ : OUTBUF
      port map(D => \apbo.prdata_c[10]\, PAD => apbo(10));
    
    \AHB_Master_Out_pad[217]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(217));
    
    \AHB_Master_Out_pad[227]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(227));
    
    \AHB_Master_Out_pad[17]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[13]\, PAD => 
        AHB_Master_Out(17));
    
    \AHB_Master_Out_pad[247]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(247));
    
    \apbo_pad[87]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(87));
    
    \apbo_pad[74]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(74));
    
    \AHB_Master_Out_pad[236]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(236));
    
    \AHB_Master_Out_pad[356]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(356));
    
    \AHB_Master_Out_pad[219]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(219));
    
    \apbo_pad[42]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(42));
    
    \AHB_Master_Out_pad[229]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(229));
    
    \AHB_Master_Out_pad[19]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[15]\, PAD => 
        AHB_Master_Out(19));
    
    \apbi_pad[71]\ : INBUF
      port map(PAD => apbi(71), Y => \apbi_c[71]\);
    
    \AHB_Master_Out_pad[53]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[6]\, PAD => 
        AHB_Master_Out(53));
    
    \AHB_Master_Out_pad[249]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(249));
    
    \AHB_Master_Out_pad[193]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(193));
    
    \AHB_Master_Out_pad[138]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(138));
    
    \apbi_pad[75]\ : INBUF
      port map(PAD => apbi(75), Y => \apbi_c[75]\);
    
    \AHB_Master_Out_pad[28]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[24]\, PAD => 
        AHB_Master_Out(28));
    
    \AHB_Master_Out_pad[91]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(91));
    
    \apbo_pad[83]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(83));
    
    \sdo_pad[6]\ : INBUF
      port map(PAD => sdo(6), Y => \sdo_c[6]\);
    
    \apbo_pad[11]\ : OUTBUF
      port map(D => \apbo.prdata_c[11]\, PAD => apbo(11));
    
    \AHB_Master_Out_pad[110]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(110));
    
    \apbo_pad[15]\ : OUTBUF
      port map(D => \apbo.prdata_c[15]\, PAD => apbo(15));
    
    \apbi_pad[24]\ : INBUF
      port map(PAD => apbi(24), Y => \apbi_c[24]\);
    
    \AHB_Master_Out_pad[267]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(267));
    
    \AHB_Master_Out_pad[120]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(120));
    
    \AHB_Master_Out_pad[140]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(140));
    
    \apbo_pad[40]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(40));
    
    \AHB_Master_Out_pad[20]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[16]\, PAD => 
        AHB_Master_Out(20));
    
    \AHB_Master_Out_pad[275]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(275));
    
    \AHB_Master_Out_pad[116]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(116));
    
    cnv_run_pad : INBUF
      port map(PAD => cnv_run, Y => cnv_run_c);
    
    \AHB_Master_Out_pad[280]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(280));
    
    \AHB_Master_Out_pad[269]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(269));
    
    \AHB_Master_Out_pad[126]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(126));
    
    \AHB_Master_Out_pad[185]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(185));
    
    \AHB_Master_Out_pad[146]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(146));
    
    \apbo_pad[128]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(128));
    
    \AHB_Master_Out_pad[333]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(333));
    
    \apbo_pad[56]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(56));
    
    \apbi_pad[49]\ : INBUF
      port map(PAD => apbi(49), Y => \apbi_c[49]\);
    
    \AHB_Master_Out_pad[64]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[17]\, PAD => 
        AHB_Master_Out(64));
    
    \AHB_Master_Out_pad[354]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(354));
    
    \AHB_Master_Out_pad[308]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(308));
    
    cnv_clk_pad : INBUF
      port map(PAD => cnv_clk, Y => cnv_clk_c);
    
    \AHB_Master_Out_pad[160]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(160));
    
    \apbo_pad[41]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(41));
    
    \apbo_pad[39]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(39));
    
    \apbi_pad[19]\ : INBUF
      port map(PAD => apbi(19), Y => \apbi_c[19]\);
    
    \AHB_Master_Out_pad[2]\ : OUTBUF
      port map(D => \AHB_Master_Out.htrans_c[0]\, PAD => 
        AHB_Master_Out(2));
    
    \apbo_pad[45]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(45));
    
    \apbi_pad[62]\ : INBUF
      port map(PAD => apbi(62), Y => \apbi_c[62]\);
    
    \AHB_Master_Out_pad[286]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(286));
    
    \apbi_pad[59]\ : INBUF
      port map(PAD => apbi(59), Y => \apbi_c[59]\);
    
    \AHB_Master_Out_pad[26]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[22]\, PAD => 
        AHB_Master_Out(26));
    
    \apbo_pad[29]\ : OUTBUF
      port map(D => \apbo.prdata_c[29]\, PAD => apbo(29));
    
    \AHB_Master_Out_pad[166]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(166));
    
    \AHB_Master_Out_pad[188]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(188));
    
    \AHB_Master_Out_pad[238]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(238));
    
    HCLK_pad : CLKBUF
      port map(PAD => HCLK, Y => HCLK_c);
    
    \AHB_Master_Out_pad[204]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(204));
    
    \AHB_Master_Out_pad[3]\ : OUTBUF
      port map(D => \AHB_Master_Out.htrans_c[1]\, PAD => 
        AHB_Master_Out(3));
    
    \AHB_Master_Out_pad[27]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[23]\, PAD => 
        AHB_Master_Out(27));
    
    \AHB_Master_Out_pad[255]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(255));
    
    \apbo_pad[69]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(69));
    
    \apbi_pad[60]\ : INBUF
      port map(PAD => apbi(60), Y => \apbi_c[60]\);
    
    \sdo_pad[2]\ : INBUF
      port map(PAD => sdo(2), Y => \sdo_c[2]\);
    
    \AHB_Master_Out_pad[34]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[30]\, PAD => 
        AHB_Master_Out(34));
    
    \AHB_Master_Out_pad[203]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(203));
    
    \AHB_Master_Out_pad[139]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(139));
    
    \AHB_Master_Out_pad[29]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[25]\, PAD => 
        AHB_Master_Out(29));
    
    \AHB_Master_Out_pad[101]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(101));
    
    \AHB_Master_Out_pad[63]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[16]\, PAD => 
        AHB_Master_Out(63));
    
    \apbo_pad[109]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(109));
    
    \apbo_pad[54]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(54));
    
    \apbo_pad[77]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(77));
    
    \apbi_pad[61]\ : INBUF
      port map(PAD => apbi(61), Y => \apbi_c[61]\);
    
    \AHB_Master_Out_pad[330]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(330));
    
    \apbo_pad[121]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(121));
    
    \apbi_pad[65]\ : INBUF
      port map(PAD => apbi(65), Y => \apbi_c[65]\);
    
    \AHB_Master_Out_pad[295]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(295));
    
    \apbo_pad[92]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(92));
    
    \AHB_Master_Out_pad[277]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(277));
    
    \AHB_Master_Out_pad[71]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[24]\, PAD => 
        AHB_Master_Out(71));
    
    \apbo_pad[73]\ : OUTBUF
      port map(D => \VCC\, PAD => apbo(73));
    
    \AHB_Master_Out_pad[81]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(81));
    
    \AHB_Master_Out_pad[279]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(279));
    
    \apbo_pad[125]\ : OUTBUF
      port map(D => \GND\, PAD => apbo(125));
    
    \AHB_Master_Out_pad[288]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(288));
    
    \AHB_Master_Out_pad[107]\ : OUTBUF
      port map(D => \GND\, PAD => AHB_Master_Out(107));
    
    \AHB_Master_Out_pad[48]\ : OUTBUF
      port map(D => \AHB_Master_Out.hwdata_c[1]\, PAD => 
        AHB_Master_Out(48));
    
    \AHB_Master_Out_pad[33]\ : OUTBUF
      port map(D => \AHB_Master_Out.haddr_c[29]\, PAD => 
        AHB_Master_Out(33));
    

end DEF_ARCH; 
