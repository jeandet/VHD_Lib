LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE lpp_lfr_management_apbreg_pkg IS
  
  CONSTANT ADDR_LFR_MANAGMENT_CONTROL          : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000000";
  CONSTANT ADDR_LFR_MANAGMENT_TIME_LOAD        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000001";
  CONSTANT ADDR_LFR_MANAGMENT_TIME_COARSE      : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000010";
  CONSTANT ADDR_LFR_MANAGMENT_TIME_FINE        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000011";
  CONSTANT ADDR_LFR_MANAGMENT_HK_TEMP_0        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000100";
  CONSTANT ADDR_LFR_MANAGMENT_HK_TEMP_1        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000101";
  CONSTANT ADDR_LFR_MANAGMENT_HK_TEMP_2        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000110";
  
END lpp_lfr_management_apbreg_pkg;
