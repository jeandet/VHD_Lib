------------------------------------------------------------------------------
--  LEON3 Demonstration design test bench
--  Copyright (C) 2004 Jiri Gaisler, Gaisler Research
------------------------------------------------------------------------------
------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2014, Aeroflex Gaisler
--  Copyright (C) 2015 - 2016, Cobham Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gaisler;
use gaisler.libdcom.all;
use gaisler.sim.all;
use work.debug.all;
library techmap;
use techmap.gencomp.all;
library micron;
use micron.components.all;
library grlib;
use grlib.stdlib.all;

use work.config.all;	-- configuration


entity testbench is
  generic (
    fabtech   : integer := CFG_FABTECH;
    memtech   : integer := CFG_MEMTECH;
    padtech   : integer := CFG_PADTECH;
    clktech   : integer := CFG_CLKTECH;
    disas     : integer := CFG_DISAS;	-- Enable disassembly to console
    dbguart   : integer := CFG_DUART;	-- Print UART on console
    pclow     : integer := CFG_PCLOW;

    clkperiod : integer := 20;		-- system clock period
    romdepth  : integer := 22		-- rom address depth (flash 4 MB)
 --   sramwidth  : integer := 32;		-- ram data width (8/16/32)
 --   sramdepth  : integer := 20;		-- ram address depth
 --   srambanks  : integer := 2		-- number of ram banks
  );
end;

architecture behav of testbench is

constant promfile  : string := "prom.srec";  -- rom contents
constant sramfile  : string := "ram.srec";  -- ram contents
constant sdramfile : string := "ram.srec"; -- sdram contents


signal SW     : std_logic_vector(4 downto 1);
signal clk : std_logic := '0';
signal Rst    : std_logic := '0';			-- Reset
constant ct : integer := clkperiod/2;

signal address  : std_logic_vector(21 downto 0);
signal data     : std_logic_vector(31 downto 24);

signal romsn    : std_logic;
signal oen      : std_logic;
signal writen   : std_logic;
signal dsuen, dsutx, dsurx, dsubre, dsuact : std_logic;
signal dsurst   : std_logic;
signal error    : std_logic;

signal sdcke    : std_logic;
signal sdcsn    : std_logic;
signal sdwen    : std_logic;                       -- write en
signal sdrasn   : std_logic;                       -- row addr stb
signal sdcasn   : std_logic;                       -- col addr stb
signal dram_ldqm : std_logic;
signal dram_udqm : std_logic;
signal sdclk    : std_logic;
signal dram_ba  : std_logic_vector(1 downto 0);

signal FTDI_RXF    :  std_logic;
signal FTDI_TXE    :  std_logic;
signal FTDI_SIWUA  :  std_logic;
signal FTDI_WR     :  std_logic;
signal FTDI_RD     :  std_logic;
signal FTDI_D      :  std_logic_vector(7 downto 0):=(others=>'Z');

constant lresp : boolean := false;


signal sa      	: std_logic_vector(12 downto 0);
signal sd   	: std_logic_vector(15 downto 0);


begin

  clk <= not clk after ct * 1 ns; --50 MHz clk
  rst <= dsurst; --reset
  dsuen <= '1';
  dsubre <= '1'; -- inverted on the board
  sw(1) <= rst;

  d3 : entity work.leon3mp
        generic map ( fabtech, memtech, padtech, clktech, disas, dbguart, pclow )
        port map (
            CLK50  => clk,
            LEDS   => open,
            SW     => SW,
            dram_addr => sa,
            dram_ba_0	=> dram_ba(0),
            dram_ba_1	=> dram_ba(1),
            dram_dq	=> sd(15 downto 0),
            dram_clk  	=> sdclk,
            dram_cke  	=> sdcke,
            dram_cs_n   => sdcsn,
            dram_we_n  	=> sdwen,
            dram_ras_n  => sdrasn,
            dram_cas_n  => sdcasn,
            dram_ldqm	  => dram_ldqm,
            dram_udqm	  => dram_udqm,
            uart_txd  	=> dsutx,
            uart_rxd  	=> dsurx,

            FTDI_RXF    => FTDI_RXF,
            FTDI_TXE    => FTDI_TXE,
            FTDI_SIWUA  => FTDI_SIWUA,
            FTDI_WR     => FTDI_WR,
            FTDI_RD     => FTDI_RD,
            FTDI_D      => FTDI_D
            );

    u1: entity work.mt48lc16m16a2 generic map (addr_bits => 13, col_bits => 9, index => 1024, fname => sdramfile)
	PORT MAP(
            Dq => sd(15 downto 0), Addr => sa(12 downto 0),
            Ba => dram_ba, Clk => sdclk, Cke => sdcke,
            Cs_n => sdcsn, Ras_n => sdrasn, Cas_n => sdcasn, We_n => sdwen,
            Dqm(0) => dram_ldqm, Dqm(1) => dram_udqm );



  error <= 'H';			  -- ERROR pull-up

   iuerr : process
   begin
     wait for 2500 ns;
     if to_x01(error) = '1' then wait on error; end if;
     assert (to_x01(error) = '1')
       report "*** IU in error mode, simulation halted ***"
         severity failure ;
   end process;

  data <= buskeep(data) after 5 ns;
  sd <= buskeep(sd) after 5 ns;

  testftdi : process
    procedure ftdi_write(signal FTDI_RXF : out std_logic; signal FTDI_RD : in std_logic;  value : integer; signal FTDI_D: out std_logic_vector(7 downto 0)) is
    begin
        FTDI_RXF <= '0';
        wait until FTDI_RD = '0';
        wait for 14 ns;
        FTDI_D <= conv_std_logic_vector(value,8);
        wait for 16 ns;
        FTDI_D <= (others=>'Z');
        wait until FTDI_RD = '1';
        FTDI_RXF <= '1';
        wait for 3 ns;
    end;
    procedure dcom_ftdi_write_reg(signal FTDI_RXF : out std_logic; signal FTDI_RD : in std_logic; address : std_logic_vector(31 downto 0); value :  std_logic_vector(31 downto 0); signal FTDI_D: out std_logic_vector(7 downto 0)) is
    begin
        ftdi_write(FTDI_RXF,FTDI_RD,16#C0#,FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(31 downto 24))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(23 downto 16))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(15 downto 8))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(7 downto 0))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(value(31 downto 24))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(value(23 downto 16))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(value(15 downto 8))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(value(7 downto 0))),FTDI_D);

    end;
    procedure dcom_ftdi_read_reg(signal FTDI_RXF : out std_logic; signal FTDI_RD : in std_logic; address : std_logic_vector(31 downto 0); signal FTDI_D: out std_logic_vector(7 downto 0)) is
    begin
        ftdi_write(FTDI_RXF,FTDI_RD,16#80#,FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(31 downto 24))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(23 downto 16))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(15 downto 8))),FTDI_D);
        ftdi_write(FTDI_RXF,FTDI_RD,to_integer(UNSIGNED(address(7 downto 0))),FTDI_D);
    end;
    begin
      FTDI_D <= (others=>'Z');
      dsurst <= '0';
      FTDI_RXF <= '1';
      wait for 100 ns;
      dsurst <= '1';
      wait for 100 ns;
      dcom_ftdi_read_reg(FTDI_RXF,FTDI_RD,X"80000000",FTDI_D);
      dcom_ftdi_read_reg(FTDI_RXF,FTDI_RD,X"80000004",FTDI_D);
      dcom_ftdi_read_reg(FTDI_RXF,FTDI_RD,X"80000008",FTDI_D);
      dcom_ftdi_read_reg(FTDI_RXF,FTDI_RD,X"8000000C",FTDI_D);
      dcom_ftdi_read_reg(FTDI_RXF,FTDI_RD,X"80000010",FTDI_D);
      wait;
 end process;

 txe: process
  begin
    FTDI_TXE <= '0';
    wait until FTDI_WR = '0';
    wait for 14 ns;
    FTDI_TXE <= '1';
    wait for 49 ns;
 end process;
end ;

