LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE lpp_lfr_apbreg_pkg IS

  -----------------------------------------------------------------------------
  -- SPECTRAL_MATRIX
  -----------------------------------------------------------------------------
  CONSTANT ADDR_LFR_SM_CONFIG           : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000000";
  CONSTANT ADDR_LFR_SM_STATUS           : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000001";
  CONSTANT ADDR_LFR_SM_F0_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000010";
  CONSTANT ADDR_LFR_SM_F0_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000011";
  
  CONSTANT ADDR_LFR_SM_F1_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000100";
  CONSTANT ADDR_LFR_SM_F1_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000101";
  CONSTANT ADDR_LFR_SM_F2_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000110";
  CONSTANT ADDR_LFR_SM_F2_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "000111";

  CONSTANT ADDR_LFR_SM_F0_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001000";
  CONSTANT ADDR_LFR_SM_F0_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001001";
  CONSTANT ADDR_LFR_SM_F0_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001010";
  CONSTANT ADDR_LFR_SM_F0_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001011";

  CONSTANT ADDR_LFR_SM_F1_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001100";
  CONSTANT ADDR_LFR_SM_F1_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001101";
  CONSTANT ADDR_LFR_SM_F1_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001110";
  CONSTANT ADDR_LFR_SM_F1_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "001111";

  CONSTANT ADDR_LFR_SM_F2_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010000";
  CONSTANT ADDR_LFR_SM_F2_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010001";
  CONSTANT ADDR_LFR_SM_F2_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010010";
  CONSTANT ADDR_LFR_SM_F2_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010011";

  CONSTANT ADDR_LFR_SM_LENGTH           : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010100";
  -----------------------------------------------------------------------------
  -- WAVEFORM PICKER
  -----------------------------------------------------------------------------
  CONSTANT ADDR_LFR_WP_DATASHAPING      : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010101";
  CONSTANT ADDR_LFR_WP_CONTROL          : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010110";
  CONSTANT ADDR_LFR_WP_F0_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "010111";

  CONSTANT ADDR_LFR_WP_F0_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011000";
  CONSTANT ADDR_LFR_WP_F1_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011001";
  CONSTANT ADDR_LFR_WP_F1_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011010";
  CONSTANT ADDR_LFR_WP_F2_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011011";

  CONSTANT ADDR_LFR_WP_F2_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011100";
  CONSTANT ADDR_LFR_WP_F3_0_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011101";
  CONSTANT ADDR_LFR_WP_F3_1_ADDR        : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011110";
  CONSTANT ADDR_LFR_WP_STATUS           : STD_LOGIC_VECTOR(7 DOWNTO 2) := "011111";

  CONSTANT ADDR_LFR_WP_DELTASNAPSHOT    : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100000";
  CONSTANT ADDR_LFR_WP_DELTA_F0         : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100001";
  CONSTANT ADDR_LFR_WP_DELTA_F0_2       : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100010";
  CONSTANT ADDR_LFR_WP_DELTA_F1         : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100011";

  CONSTANT ADDR_LFR_WP_DELTA_F2         : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100100";
  CONSTANT ADDR_LFR_WP_DATA_IN_BUFFER   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100101";
  CONSTANT ADDR_LFR_WP_NBSNAPSHOT       : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100110";
  CONSTANT ADDR_LFR_WP_START_DATE       : STD_LOGIC_VECTOR(7 DOWNTO 2) := "100111";

  CONSTANT ADDR_LFR_WP_F0_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101000";
  CONSTANT ADDR_LFR_WP_F0_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101001";
  CONSTANT ADDR_LFR_WP_F0_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101010";
  CONSTANT ADDR_LFR_WP_F0_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101011";

  CONSTANT ADDR_LFR_WP_F1_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101100";
  CONSTANT ADDR_LFR_WP_F1_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101101";
  CONSTANT ADDR_LFR_WP_F1_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101110";
  CONSTANT ADDR_LFR_WP_F1_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "101111";

  CONSTANT ADDR_LFR_WP_F2_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110000";
  CONSTANT ADDR_LFR_WP_F2_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110001";
  CONSTANT ADDR_LFR_WP_F2_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110010";
  CONSTANT ADDR_LFR_WP_F2_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110011";

  CONSTANT ADDR_LFR_WP_F3_0_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110100";
  CONSTANT ADDR_LFR_WP_F3_0_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110101";
  CONSTANT ADDR_LFR_WP_F3_1_TIME_COARSE : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110110";
  CONSTANT ADDR_LFR_WP_F3_1_TIME_FINE   : STD_LOGIC_VECTOR(7 DOWNTO 2) := "110111";

  CONSTANT ADDR_LFR_WP_LENGTH           : STD_LOGIC_VECTOR(7 DOWNTO 2) := "111000";  
  -----------------------------------------------------------------------------
  -- LFR
  -----------------------------------------------------------------------------
  CONSTANT ADDR_LFR_VERSION             : STD_LOGIC_VECTOR(7 DOWNTO 2) := "111100";  
  

END lpp_lfr_apbreg_pkg;
